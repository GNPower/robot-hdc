`timescale 1ns/100ps

module Bundler
(
	// clock and reset
	clk,
	reset_n,
	
	// Input data
	start,
	
	// Output data
	done
);


endmodule
