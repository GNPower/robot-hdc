module fp_accum (
		input  wire        clk,    //    clk.clk
		input  wire        areset, // areset.reset
		input  wire [31:0] a,      //      a.a
		output wire [31:0] q,      //      q.q
		input  wire [0:0]  acc     //    acc.acc
	);
endmodule

