// Copyright (C) 2019  Intel Corporation. All rights reserved.
// Your use of Intel Corporation's design tools, logic functions 
// and other software and tools, and any partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Intel Program License 
// Subscription Agreement, the Intel Quartus Prime License Agreement,
// the Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is for
// the sole purpose of programming logic devices manufactured by
// Intel and sold by Intel or its authorized distributors.  Please
// refer to the applicable agreement for further details, at
// https://fpgasoftware.intel.com/eula.

// VENDOR "Altera"
// PROGRAM "Quartus Prime"
// VERSION "Version 19.1.0 Build 240 03/26/2019 SJ Pro Edition"

// DATE "11/01/2023 17:17:25"

// 
// Device: Altera 1SG280HN1F43E2VGS1 Package FBGA1760
// 

// 
// This greybox netlist file is for third party Synthesis Tools
// for timing and resource estimation only.
// 


module fp_add (
	q,
	clk,
	areset,
	b,
	a)/* synthesis synthesis_greybox=0 */;
output 	[31:0] q;
input 	clk;
input 	areset;
input 	[31:0] b;
input 	[31:0] a;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire fp_functions_0_aredist2_aMinusA_uid87_fpAddTest_q_1_q_a0_a_aq;
wire fp_functions_0_aregInputs_uid118_fpAddTest_delay_adelay_signals_a0_a_a0_a_aq;
wire fp_functions_0_aredist16_excZ_aSig_uid16_uid23_fpAddTest_q_1_q_a0_a_aq;
wire fp_functions_0_aredist14_excZ_bSig_uid17_uid37_fpAddTest_q_3_q_a0_a_aq;
wire fp_functions_0_aredist4_effSub_uid52_fpAddTest_q_2_q_a0_a_aq;
wire fp_functions_0_aredist15_excI_aSig_uid27_fpAddTest_q_1_q_a0_a_aq;
wire fp_functions_0_aredist10_excI_bSig_uid41_fpAddTest_q_1_q_a0_a_aq;
wire fp_functions_0_aexcN_bSig_uid42_fpAddTest_delay_adelay_signals_a0_a_a0_a_aq;
wire fp_functions_0_aexcN_aSig_uid28_fpAddTest_delay_adelay_signals_a0_a_a0_a_aq;
wire fp_functions_0_aadd_7_a1_sumout;
wire fp_functions_0_aadd_7_a2;
wire fp_functions_0_aadd_7_a6_sumout;
wire fp_functions_0_aadd_7_a7;
wire fp_functions_0_aadd_7_a11_sumout;
wire fp_functions_0_aadd_7_a12;
wire fp_functions_0_aadd_7_a16_sumout;
wire fp_functions_0_aadd_7_a17;
wire fp_functions_0_aadd_7_a21_sumout;
wire fp_functions_0_aadd_7_a22;
wire fp_functions_0_aadd_7_a26_sumout;
wire fp_functions_0_aadd_7_a27;
wire fp_functions_0_aadd_7_a31_sumout;
wire fp_functions_0_aadd_7_a32;
wire fp_functions_0_aadd_7_a36_sumout;
wire fp_functions_0_aadd_7_a37;
wire fp_functions_0_aadd_7_a41_sumout;
wire fp_functions_0_aadd_7_a42;
wire fp_functions_0_aadd_7_a46_sumout;
wire fp_functions_0_aadd_7_a47;
wire fp_functions_0_aadd_7_a51_sumout;
wire fp_functions_0_aadd_7_a56_sumout;
wire fp_functions_0_aadd_7_a57;
wire fp_functions_0_aadd_7_a61_sumout;
wire fp_functions_0_aadd_7_a62;
wire fp_functions_0_aadd_7_a66_sumout;
wire fp_functions_0_aadd_7_a67;
wire fp_functions_0_aadd_7_a71_sumout;
wire fp_functions_0_aadd_7_a72;
wire fp_functions_0_aadd_7_a76_sumout;
wire fp_functions_0_aadd_7_a77;
wire fp_functions_0_aadd_7_a81_sumout;
wire fp_functions_0_aadd_7_a82;
wire fp_functions_0_aadd_7_a86_sumout;
wire fp_functions_0_aadd_7_a87;
wire fp_functions_0_aadd_7_a91_sumout;
wire fp_functions_0_aadd_7_a92;
wire fp_functions_0_aadd_7_a96_sumout;
wire fp_functions_0_aadd_7_a97;
wire fp_functions_0_aadd_7_a101_sumout;
wire fp_functions_0_aadd_7_a102;
wire fp_functions_0_aadd_7_a106_sumout;
wire fp_functions_0_aadd_7_a107;
wire fp_functions_0_aadd_7_a111_sumout;
wire fp_functions_0_aadd_7_a112;
wire fp_functions_0_aadd_7_a116_sumout;
wire fp_functions_0_aadd_7_a117;
wire fp_functions_0_aadd_7_a121_sumout;
wire fp_functions_0_aadd_7_a122;
wire fp_functions_0_aadd_7_a126_sumout;
wire fp_functions_0_aadd_7_a127;
wire fp_functions_0_aadd_7_a131_sumout;
wire fp_functions_0_aadd_7_a132;
wire fp_functions_0_aadd_7_a136_sumout;
wire fp_functions_0_aadd_7_a137;
wire fp_functions_0_aadd_7_a141_sumout;
wire fp_functions_0_aadd_7_a142;
wire fp_functions_0_aadd_7_a146_sumout;
wire fp_functions_0_aadd_7_a147;
wire fp_functions_0_aadd_7_a151_sumout;
wire fp_functions_0_aadd_7_a152;
wire fp_functions_0_aadd_7_a156_sumout;
wire fp_functions_0_aadd_7_a157;
wire fp_functions_0_aadd_7_a161_sumout;
wire fp_functions_0_aadd_7_a162;
wire fp_functions_0_asignRInfRZRReg_uid137_fpAddTest_delay_adelay_signals_a0_a_a0_a_aq;
wire fp_functions_0_aredist1_vCount_uid152_lzCountVal_uid85_fpAddTest_q_1_q_a0_a_aq;
wire fp_functions_0_avStagei_uid157_lzCountVal_uid85_fpAddTest_q_a11_a_aq;
wire fp_functions_0_avStagei_uid157_lzCountVal_uid85_fpAddTest_q_a10_a_aq;
wire fp_functions_0_avStagei_uid157_lzCountVal_uid85_fpAddTest_q_a8_a_aq;
wire fp_functions_0_avStagei_uid157_lzCountVal_uid85_fpAddTest_q_a9_a_aq;
wire fp_functions_0_avStagei_uid157_lzCountVal_uid85_fpAddTest_q_a15_a_aq;
wire fp_functions_0_avStagei_uid157_lzCountVal_uid85_fpAddTest_q_a14_a_aq;
wire fp_functions_0_avStagei_uid157_lzCountVal_uid85_fpAddTest_q_a7_a_aq;
wire fp_functions_0_avStagei_uid157_lzCountVal_uid85_fpAddTest_q_a12_a_aq;
wire fp_functions_0_avStagei_uid157_lzCountVal_uid85_fpAddTest_q_a13_a_aq;
wire fp_functions_0_avStagei_uid157_lzCountVal_uid85_fpAddTest_q_a6_a_aq;
wire fp_functions_0_avStagei_uid157_lzCountVal_uid85_fpAddTest_q_a5_a_aq;
wire fp_functions_0_avStagei_uid157_lzCountVal_uid85_fpAddTest_q_a4_a_aq;
wire fp_functions_0_avStagei_uid157_lzCountVal_uid85_fpAddTest_q_a3_a_aq;
wire fp_functions_0_avStagei_uid157_lzCountVal_uid85_fpAddTest_q_a2_a_aq;
wire fp_functions_0_avStagei_uid157_lzCountVal_uid85_fpAddTest_q_a1_a_aq;
wire fp_functions_0_aredist12_expXIsMax_uid38_fpAddTest_q_2_q_a0_a_aq;
wire fp_functions_0_aredist9_InvExpXIsZero_uid44_fpAddTest_q_2_q_a0_a_aq;
wire fp_functions_0_aredist18_exp_aSig_uid21_fpAddTest_b_2_q_a4_a_aq;
wire fp_functions_0_aredist18_exp_aSig_uid21_fpAddTest_b_2_q_a5_a_aq;
wire fp_functions_0_aredist18_exp_aSig_uid21_fpAddTest_b_2_q_a6_a_aq;
wire fp_functions_0_aredist18_exp_aSig_uid21_fpAddTest_b_2_q_a7_a_aq;
wire fp_functions_0_aredist18_exp_aSig_uid21_fpAddTest_b_2_q_a0_a_aq;
wire fp_functions_0_aredist18_exp_aSig_uid21_fpAddTest_b_2_q_a1_a_aq;
wire fp_functions_0_aredist18_exp_aSig_uid21_fpAddTest_b_2_q_a2_a_aq;
wire fp_functions_0_aredist18_exp_aSig_uid21_fpAddTest_b_2_q_a3_a_aq;
wire fp_functions_0_aredist13_excZ_bSig_uid17_uid37_fpAddTest_q_2_q_a0_a_aq;
wire fp_functions_0_aredist4_effSub_uid52_fpAddTest_q_2_delay_0_a0_a_aq;
wire fp_functions_0_afracXIsZero_uid25_fpAddTest_delay_adelay_signals_a0_a_a0_a_aq;
wire fp_functions_0_aredist11_fracXIsZero_uid39_fpAddTest_q_2_q_a0_a_aq;
wire fp_functions_0_aleftShiftStage2_uid249_fracPostNormExt_uid88_fpAddTest_q_a4_a_aq;
wire fp_functions_0_aadd_7_a167_cout;
wire fp_functions_0_aexpPostNorm_uid92_fpAddTest_o_a5_a_aq;
wire fp_functions_0_aexpPostNorm_uid92_fpAddTest_o_a0_a_aq;
wire fp_functions_0_aexpPostNorm_uid92_fpAddTest_o_a1_a_aq;
wire fp_functions_0_aexpPostNorm_uid92_fpAddTest_o_a2_a_aq;
wire fp_functions_0_aexpPostNorm_uid92_fpAddTest_o_a3_a_aq;
wire fp_functions_0_aexpPostNorm_uid92_fpAddTest_o_a4_a_aq;
wire fp_functions_0_aexpPostNorm_uid92_fpAddTest_o_a6_a_aq;
wire fp_functions_0_aexpPostNorm_uid92_fpAddTest_o_a7_a_aq;
wire fp_functions_0_aexpPostNorm_uid92_fpAddTest_o_a8_a_aq;
wire fp_functions_0_aexpPostNorm_uid92_fpAddTest_o_a9_a_aq;
wire fp_functions_0_aleftShiftStage2_uid249_fracPostNormExt_uid88_fpAddTest_q_a5_a_aq;
wire fp_functions_0_aleftShiftStage2_uid249_fracPostNormExt_uid88_fpAddTest_q_a6_a_aq;
wire fp_functions_0_aleftShiftStage2_uid249_fracPostNormExt_uid88_fpAddTest_q_a7_a_aq;
wire fp_functions_0_aleftShiftStage2_uid249_fracPostNormExt_uid88_fpAddTest_q_a8_a_aq;
wire fp_functions_0_aleftShiftStage2_uid249_fracPostNormExt_uid88_fpAddTest_q_a9_a_aq;
wire fp_functions_0_aleftShiftStage2_uid249_fracPostNormExt_uid88_fpAddTest_q_a10_a_aq;
wire fp_functions_0_aleftShiftStage2_uid249_fracPostNormExt_uid88_fpAddTest_q_a11_a_aq;
wire fp_functions_0_aleftShiftStage2_uid249_fracPostNormExt_uid88_fpAddTest_q_a12_a_aq;
wire fp_functions_0_aleftShiftStage2_uid249_fracPostNormExt_uid88_fpAddTest_q_a13_a_aq;
wire fp_functions_0_aleftShiftStage2_uid249_fracPostNormExt_uid88_fpAddTest_q_a14_a_aq;
wire fp_functions_0_aleftShiftStage2_uid249_fracPostNormExt_uid88_fpAddTest_q_a15_a_aq;
wire fp_functions_0_aleftShiftStage2_uid249_fracPostNormExt_uid88_fpAddTest_q_a16_a_aq;
wire fp_functions_0_aleftShiftStage2_uid249_fracPostNormExt_uid88_fpAddTest_q_a17_a_aq;
wire fp_functions_0_aleftShiftStage2_uid249_fracPostNormExt_uid88_fpAddTest_q_a18_a_aq;
wire fp_functions_0_aleftShiftStage2_uid249_fracPostNormExt_uid88_fpAddTest_q_a19_a_aq;
wire fp_functions_0_aleftShiftStage2_uid249_fracPostNormExt_uid88_fpAddTest_q_a20_a_aq;
wire fp_functions_0_aleftShiftStage2_uid249_fracPostNormExt_uid88_fpAddTest_q_a21_a_aq;
wire fp_functions_0_aleftShiftStage2_uid249_fracPostNormExt_uid88_fpAddTest_q_a22_a_aq;
wire fp_functions_0_aleftShiftStage2_uid249_fracPostNormExt_uid88_fpAddTest_q_a23_a_aq;
wire fp_functions_0_aleftShiftStage2_uid249_fracPostNormExt_uid88_fpAddTest_q_a24_a_aq;
wire fp_functions_0_aleftShiftStage2_uid249_fracPostNormExt_uid88_fpAddTest_q_a25_a_aq;
wire fp_functions_0_aleftShiftStage2_uid249_fracPostNormExt_uid88_fpAddTest_q_a26_a_aq;
wire fp_functions_0_aredist6_sigB_uid51_fpAddTest_b_2_q_a0_a_aq;
wire fp_functions_0_aredist8_sigA_uid50_fpAddTest_b_2_q_a0_a_aq;
wire fp_functions_0_aadd_4_a1_sumout;
wire fp_functions_0_aadd_4_a2;
wire fp_functions_0_aadd_4_a6_sumout;
wire fp_functions_0_aadd_4_a7;
wire fp_functions_0_aadd_4_a11_sumout;
wire fp_functions_0_aadd_4_a12;
wire fp_functions_0_aadd_4_a16_sumout;
wire fp_functions_0_aadd_4_a17;
wire fp_functions_0_aadd_4_a21_sumout;
wire fp_functions_0_aadd_4_a22;
wire fp_functions_0_aadd_4_a26_sumout;
wire fp_functions_0_aadd_4_a27;
wire fp_functions_0_aadd_4_a31_sumout;
wire fp_functions_0_aadd_4_a32;
wire fp_functions_0_aadd_4_a36_sumout;
wire fp_functions_0_aadd_4_a37;
wire fp_functions_0_aadd_4_a41_sumout;
wire fp_functions_0_aadd_4_a42;
wire fp_functions_0_aadd_4_a46_sumout;
wire fp_functions_0_aadd_4_a47;
wire fp_functions_0_aadd_4_a51_sumout;
wire fp_functions_0_aadd_4_a52;
wire fp_functions_0_aadd_4_a56_sumout;
wire fp_functions_0_aadd_4_a57;
wire fp_functions_0_aadd_4_a61_sumout;
wire fp_functions_0_aadd_4_a62;
wire fp_functions_0_aadd_4_a66_sumout;
wire fp_functions_0_aadd_4_a67;
wire fp_functions_0_aadd_4_a71_sumout;
wire fp_functions_0_aadd_4_a72;
wire fp_functions_0_aadd_4_a76_sumout;
wire fp_functions_0_aadd_4_a81_sumout;
wire fp_functions_0_aadd_4_a82;
wire fp_functions_0_aadd_4_a86_sumout;
wire fp_functions_0_aadd_4_a87;
wire fp_functions_0_aadd_4_a91_sumout;
wire fp_functions_0_aadd_4_a92;
wire fp_functions_0_aadd_4_a96_sumout;
wire fp_functions_0_aadd_4_a97;
wire fp_functions_0_aadd_4_a101_sumout;
wire fp_functions_0_aadd_4_a102;
wire fp_functions_0_aadd_4_a106_sumout;
wire fp_functions_0_aadd_4_a107;
wire fp_functions_0_aadd_4_a111_sumout;
wire fp_functions_0_aadd_4_a112;
wire fp_functions_0_aadd_4_a116_sumout;
wire fp_functions_0_aadd_4_a117;
wire fp_functions_0_aadd_4_a121_sumout;
wire fp_functions_0_aadd_4_a122;
wire fp_functions_0_aadd_4_a126_sumout;
wire fp_functions_0_aadd_4_a127;
wire fp_functions_0_aadd_4_a131_sumout;
wire fp_functions_0_aadd_4_a132;
wire fp_functions_0_ashiftedOut_uid63_fpAddTest_o_a10_a_aq;
wire fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a22_a_aq;
wire fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a16_a_aq;
wire fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a0_a_aq;
wire fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a1_a_aq;
wire fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a9_a_aq;
wire fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a4_a_aq;
wire fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a21_a_aq;
wire fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a20_a_aq;
wire fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a19_a_aq;
wire fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a17_a_aq;
wire fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a18_a_aq;
wire fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a8_a_aq;
wire fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a7_a_aq;
wire fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a6_a_aq;
wire fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a5_a_aq;
wire fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a2_a_aq;
wire fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a3_a_aq;
wire fp_functions_0_aexpXIsMax_uid38_fpAddTest_delay_adelay_signals_a0_a_a0_a_aq;
wire fp_functions_0_aredist9_InvExpXIsZero_uid44_fpAddTest_q_2_delay_0_a0_a_aq;
wire fp_functions_0_aredist18_exp_aSig_uid21_fpAddTest_b_2_delay_0_a4_a_aq;
wire fp_functions_0_aredist18_exp_aSig_uid21_fpAddTest_b_2_delay_0_a5_a_aq;
wire fp_functions_0_aredist18_exp_aSig_uid21_fpAddTest_b_2_delay_0_a6_a_aq;
wire fp_functions_0_aredist18_exp_aSig_uid21_fpAddTest_b_2_delay_0_a7_a_aq;
wire fp_functions_0_aredist18_exp_aSig_uid21_fpAddTest_b_2_delay_0_a0_a_aq;
wire fp_functions_0_aredist18_exp_aSig_uid21_fpAddTest_b_2_delay_0_a1_a_aq;
wire fp_functions_0_aredist18_exp_aSig_uid21_fpAddTest_b_2_delay_0_a2_a_aq;
wire fp_functions_0_aredist18_exp_aSig_uid21_fpAddTest_b_2_delay_0_a3_a_aq;
wire fp_functions_0_aredist13_excZ_bSig_uid17_uid37_fpAddTest_q_2_delay_0_a0_a_aq;
wire fp_functions_0_aredist7_sigA_uid50_fpAddTest_b_1_q_a0_a_aq;
wire fp_functions_0_aredist5_sigB_uid51_fpAddTest_b_1_q_a0_a_aq;
wire fp_functions_0_aredist17_frac_aSig_uid22_fpAddTest_b_1_q_a19_a_aq;
wire fp_functions_0_aredist17_frac_aSig_uid22_fpAddTest_b_1_q_a21_a_aq;
wire fp_functions_0_aredist17_frac_aSig_uid22_fpAddTest_b_1_q_a15_a_aq;
wire fp_functions_0_aredist17_frac_aSig_uid22_fpAddTest_b_1_q_a16_a_aq;
wire fp_functions_0_aredist17_frac_aSig_uid22_fpAddTest_b_1_q_a17_a_aq;
wire fp_functions_0_aredist17_frac_aSig_uid22_fpAddTest_b_1_q_a18_a_aq;
wire fp_functions_0_aredist17_frac_aSig_uid22_fpAddTest_b_1_q_a20_a_aq;
wire fp_functions_0_aredist17_frac_aSig_uid22_fpAddTest_b_1_q_a22_a_aq;
wire fp_functions_0_aredist17_frac_aSig_uid22_fpAddTest_b_1_q_a2_a_aq;
wire fp_functions_0_aredist17_frac_aSig_uid22_fpAddTest_b_1_q_a0_a_aq;
wire fp_functions_0_aredist17_frac_aSig_uid22_fpAddTest_b_1_q_a1_a_aq;
wire fp_functions_0_aredist17_frac_aSig_uid22_fpAddTest_b_1_q_a8_a_aq;
wire fp_functions_0_aredist17_frac_aSig_uid22_fpAddTest_b_1_q_a13_a_aq;
wire fp_functions_0_aredist17_frac_aSig_uid22_fpAddTest_b_1_q_a14_a_aq;
wire fp_functions_0_aredist17_frac_aSig_uid22_fpAddTest_b_1_q_a9_a_aq;
wire fp_functions_0_aredist17_frac_aSig_uid22_fpAddTest_b_1_q_a10_a_aq;
wire fp_functions_0_aredist17_frac_aSig_uid22_fpAddTest_b_1_q_a11_a_aq;
wire fp_functions_0_aredist17_frac_aSig_uid22_fpAddTest_b_1_q_a12_a_aq;
wire fp_functions_0_aredist17_frac_aSig_uid22_fpAddTest_b_1_q_a3_a_aq;
wire fp_functions_0_aredist17_frac_aSig_uid22_fpAddTest_b_1_q_a4_a_aq;
wire fp_functions_0_aredist17_frac_aSig_uid22_fpAddTest_b_1_q_a5_a_aq;
wire fp_functions_0_aredist17_frac_aSig_uid22_fpAddTest_b_1_q_a6_a_aq;
wire fp_functions_0_aredist17_frac_aSig_uid22_fpAddTest_b_1_q_a7_a_aq;
wire fp_functions_0_afracXIsZero_uid39_fpAddTest_delay_adelay_signals_a0_a_a0_a_aq;
wire fp_functions_0_aredist0_vStage_uid154_lzCountVal_uid85_fpAddTest_b_1_q_a0_a_aq;
wire fp_functions_0_aredist0_vStage_uid154_lzCountVal_uid85_fpAddTest_b_1_q_a3_a_aq;
wire fp_functions_0_aredist0_vStage_uid154_lzCountVal_uid85_fpAddTest_b_1_q_a1_a_aq;
wire fp_functions_0_aredist0_vStage_uid154_lzCountVal_uid85_fpAddTest_b_1_q_a4_a_aq;
wire fp_functions_0_aredist0_vStage_uid154_lzCountVal_uid85_fpAddTest_b_1_q_a2_a_aq;
wire fp_functions_0_aleftShiftStage2_uid249_fracPostNormExt_uid88_fpAddTest_q_a3_a_aq;
wire fp_functions_0_aleftShiftStage2_uid249_fracPostNormExt_uid88_fpAddTest_q_a2_a_aq;
wire fp_functions_0_aleftShiftStage2_uid249_fracPostNormExt_uid88_fpAddTest_q_a0_a_aq;
wire fp_functions_0_aleftShiftStage2_uid249_fracPostNormExt_uid88_fpAddTest_q_a1_a_aq;
wire fp_functions_0_aadd_6_a1_sumout;
wire fp_functions_0_aadd_6_a2;
wire fp_functions_0_aadd_6_a6_sumout;
wire fp_functions_0_aadd_6_a7;
wire fp_functions_0_aadd_6_a11_sumout;
wire fp_functions_0_aadd_6_a12;
wire fp_functions_0_aadd_6_a16_sumout;
wire fp_functions_0_aadd_6_a17;
wire fp_functions_0_aadd_6_a21_sumout;
wire fp_functions_0_aadd_6_a22;
wire fp_functions_0_aadd_6_a26_sumout;
wire fp_functions_0_aadd_6_a27;
wire fp_functions_0_aadd_6_a31_sumout;
wire fp_functions_0_aadd_6_a32;
wire fp_functions_0_aadd_6_a36_sumout;
wire fp_functions_0_aadd_6_a37;
wire fp_functions_0_aadd_6_a41_sumout;
wire fp_functions_0_aadd_6_a42;
wire fp_functions_0_aadd_6_a46_sumout;
wire fp_functions_0_aredist0_vStage_uid154_lzCountVal_uid85_fpAddTest_b_1_q_a5_a_aq;
wire fp_functions_0_aredist0_vStage_uid154_lzCountVal_uid85_fpAddTest_b_1_q_a6_a_aq;
wire fp_functions_0_aredist0_vStage_uid154_lzCountVal_uid85_fpAddTest_b_1_q_a7_a_aq;
wire fp_functions_0_aredist0_vStage_uid154_lzCountVal_uid85_fpAddTest_b_1_q_a8_a_aq;
wire fp_functions_0_aredist0_vStage_uid154_lzCountVal_uid85_fpAddTest_b_1_q_a9_a_aq;
wire fp_functions_0_aredist0_vStage_uid154_lzCountVal_uid85_fpAddTest_b_1_q_a10_a_aq;
wire fp_functions_0_aredist3_fracGRS_uid84_fpAddTest_q_1_q_a11_a_aq;
wire fp_functions_0_aredist3_fracGRS_uid84_fpAddTest_q_1_q_a12_a_aq;
wire fp_functions_0_aredist3_fracGRS_uid84_fpAddTest_q_1_q_a13_a_aq;
wire fp_functions_0_aredist3_fracGRS_uid84_fpAddTest_q_1_q_a14_a_aq;
wire fp_functions_0_aredist3_fracGRS_uid84_fpAddTest_q_1_q_a15_a_aq;
wire fp_functions_0_aredist3_fracGRS_uid84_fpAddTest_q_1_q_a16_a_aq;
wire fp_functions_0_aredist3_fracGRS_uid84_fpAddTest_q_1_q_a17_a_aq;
wire fp_functions_0_aredist3_fracGRS_uid84_fpAddTest_q_1_q_a18_a_aq;
wire fp_functions_0_aredist3_fracGRS_uid84_fpAddTest_q_1_q_a19_a_aq;
wire fp_functions_0_aredist3_fracGRS_uid84_fpAddTest_q_1_q_a20_a_aq;
wire fp_functions_0_aredist3_fracGRS_uid84_fpAddTest_q_1_q_a21_a_aq;
wire fp_functions_0_aredist3_fracGRS_uid84_fpAddTest_q_1_q_a22_a_aq;
wire fp_functions_0_aredist3_fracGRS_uid84_fpAddTest_q_1_q_a23_a_aq;
wire fp_functions_0_aredist3_fracGRS_uid84_fpAddTest_q_1_q_a24_a_aq;
wire fp_functions_0_aredist3_fracGRS_uid84_fpAddTest_q_1_q_a25_a_aq;
wire fp_functions_0_aredist3_fracGRS_uid84_fpAddTest_q_1_q_a26_a_aq;
wire fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a42_a_aq;
wire fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a38_a_aq;
wire fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a34_a_aq;
wire fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a35_a_aq;
wire fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a36_a_aq;
wire fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a37_a_aq;
wire fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a39_a_aq;
wire fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a40_a_aq;
wire fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a41_a_aq;
wire fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a47_a_aq;
wire fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a48_a_aq;
wire fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a43_a_aq;
wire fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a44_a_aq;
wire fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a45_a_aq;
wire fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a46_a_aq;
wire fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a29_a_aq;
wire fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a28_a_aq;
wire fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a26_a_aq;
wire fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a27_a_aq;
wire fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a33_a_aq;
wire fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a32_a_aq;
wire fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a25_a_aq;
wire fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a30_a_aq;
wire fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a31_a_aq;
wire fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a24_a_aq;
wire fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a23_a_aq;
wire fp_functions_0_aadd_2_a1_sumout;
wire fp_functions_0_aadd_1_a1_sumout;
wire fp_functions_0_aadd_1_a2;
wire fp_functions_0_aadd_1_a6_sumout;
wire fp_functions_0_aadd_1_a7;
wire fp_functions_0_aadd_1_a11_sumout;
wire fp_functions_0_aadd_1_a12;
wire fp_functions_0_aadd_0_a1_sumout;
wire fp_functions_0_aadd_1_a16_sumout;
wire fp_functions_0_aadd_1_a17;
wire fp_functions_0_aadd_1_a21_sumout;
wire fp_functions_0_aadd_1_a22;
wire fp_functions_0_aadd_1_a26_sumout;
wire fp_functions_0_aadd_1_a27;
wire fp_functions_0_aadd_3_a1_sumout;
wire fp_functions_0_aadd_5_a1_sumout;
wire fp_functions_0_aadd_5_a2;
wire fp_functions_0_aadd_5_a6_sumout;
wire fp_functions_0_aadd_5_a7;
wire fp_functions_0_aadd_6_a52_cout;
wire fp_functions_0_aadd_5_a11_sumout;
wire fp_functions_0_aadd_5_a12;
wire fp_functions_0_aadd_5_a16_sumout;
wire fp_functions_0_aadd_5_a17;
wire fp_functions_0_aadd_5_a21_sumout;
wire fp_functions_0_aadd_5_a22;
wire fp_functions_0_aadd_5_a26_sumout;
wire fp_functions_0_aadd_5_a27;
wire fp_functions_0_aadd_5_a31_sumout;
wire fp_functions_0_aadd_5_a32;
wire fp_functions_0_aadd_5_a36_sumout;
wire fp_functions_0_aadd_5_a37;
wire fp_functions_0_aadd_5_a41_sumout;
wire fp_functions_0_aadd_2_a7_cout;
wire fp_functions_0_aadd_1_a32_cout;
wire fp_functions_0_aadd_0_a7_cout;
wire fp_functions_0_aadd_3_a7_cout;
wire fp_functions_0_aadd_1_a36_sumout;
wire fp_functions_0_aadd_2_a12_cout;
wire fp_functions_0_aadd_0_a12_cout;
wire fp_functions_0_aadd_3_a12_cout;
wire fp_functions_0_aadd_1_a41_sumout;
wire fp_functions_0_aadd_1_a42;
wire fp_functions_0_aadd_2_a17_cout;
wire fp_functions_0_aadd_0_a17_cout;
wire fp_functions_0_aadd_3_a17_cout;
wire fp_functions_0_aadd_1_a46_sumout;
wire fp_functions_0_aadd_1_a47;
wire fp_functions_0_aadd_2_a22_cout;
wire fp_functions_0_aadd_0_a22_cout;
wire fp_functions_0_aadd_3_a22_cout;
wire fp_functions_0_aadd_2_a27_cout;
wire fp_functions_0_aadd_0_a27_cout;
wire fp_functions_0_aadd_3_a27_cout;
wire fp_functions_0_aadd_2_a32_cout;
wire fp_functions_0_aadd_0_a32_cout;
wire fp_functions_0_aadd_3_a32_cout;
wire fp_functions_0_aadd_2_a37_cout;
wire fp_functions_0_aadd_0_a37_cout;
wire fp_functions_0_aadd_3_a37_cout;
wire fp_functions_0_aadd_2_a42_cout;
wire fp_functions_0_aadd_0_a42_cout;
wire fp_functions_0_aadd_3_a42_cout;
wire fp_functions_0_aadd_2_a47_cout;
wire fp_functions_0_aadd_0_a47_cout;
wire fp_functions_0_aadd_3_a47_cout;
wire fp_functions_0_aadd_2_a52_cout;
wire fp_functions_0_aadd_0_a52_cout;
wire fp_functions_0_aadd_0_a57_cout;
wire fp_functions_0_aadd_0_a62_cout;
wire fp_functions_0_aadd_0_a67_cout;
wire fp_functions_0_aadd_0_a72_cout;
wire fp_functions_0_aadd_0_a77_cout;
wire fp_functions_0_aadd_0_a82_cout;
wire fp_functions_0_aadd_0_a87_cout;
wire fp_functions_0_aadd_0_a92_cout;
wire fp_functions_0_aadd_0_a97_cout;
wire fp_functions_0_aadd_0_a102_cout;
wire fp_functions_0_aadd_0_a107_cout;
wire fp_functions_0_aadd_0_a112_cout;
wire fp_functions_0_aadd_0_a117_cout;
wire fp_functions_0_aadd_0_a122_cout;
wire fp_functions_0_aadd_0_a127_cout;
wire fp_functions_0_aadd_0_a132_cout;
wire fp_functions_0_aadd_0_a137_cout;
wire fp_functions_0_aadd_0_a142_cout;
wire fp_functions_0_aadd_0_a147_cout;
wire fp_functions_0_aadd_0_a152_cout;
wire fp_functions_0_aadd_0_a157_cout;
wire fp_functions_0_aadd_0_a162_cout;
wire fp_functions_0_areduce_nor_7_a3_combout;
wire fp_functions_0_ai1783_a34_combout;
wire fp_functions_0_ai1783_a39_combout;
wire fp_functions_0_aMux_55_a1_combout;
wire fp_functions_0_ai1783_a44_combout;
wire fp_functions_0_ai1783_a49_combout;
wire fp_functions_0_aMux_204_a0_combout;
wire fp_functions_0_aMux_236_a0_combout;
wire fp_functions_0_areduce_nor_15_a0_combout;
wire fp_functions_0_aexcRZeroVInC_uid119_fpAddTest_q_a3_a_acombout;
wire fp_functions_0_aMux_204_a1_combout;
wire fp_functions_0_aexcRInfVInC_uid122_fpAddTest_q_a5_a_a0_combout;
wire fp_functions_0_aexcRInfVInC_uid122_fpAddTest_q_a5_a_a1_combout;
wire fp_functions_0_aMux_203_a2_combout;
wire fp_functions_0_aMux_237_a2_combout;
wire fp_functions_0_aMux_236_a1_combout;
wire fp_functions_0_aMux_235_a0_combout;
wire fp_functions_0_aMux_234_a0_combout;
wire fp_functions_0_aMux_233_a0_combout;
wire fp_functions_0_aMux_232_a0_combout;
wire fp_functions_0_aMux_231_a0_combout;
wire fp_functions_0_aMux_230_a0_combout;
wire fp_functions_0_aMux_229_a0_combout;
wire fp_functions_0_aMux_228_a0_combout;
wire fp_functions_0_aMux_227_a0_combout;
wire fp_functions_0_aMux_226_a0_combout;
wire fp_functions_0_aMux_225_a0_combout;
wire fp_functions_0_aMux_224_a0_combout;
wire fp_functions_0_aMux_223_a0_combout;
wire fp_functions_0_aMux_222_a0_combout;
wire fp_functions_0_aMux_221_a0_combout;
wire fp_functions_0_aMux_220_a0_combout;
wire fp_functions_0_aMux_219_a0_combout;
wire fp_functions_0_aMux_218_a0_combout;
wire fp_functions_0_aMux_217_a0_combout;
wire fp_functions_0_aMux_216_a0_combout;
wire fp_functions_0_aMux_215_a0_combout;
wire fp_functions_0_aMux_214_a2_combout;
wire fp_functions_0_aMux_213_a2_combout;
wire fp_functions_0_aMux_212_a2_combout;
wire fp_functions_0_aMux_211_a2_combout;
wire fp_functions_0_aMux_210_a2_combout;
wire fp_functions_0_aMux_209_a2_combout;
wire fp_functions_0_aMux_208_a2_combout;
wire fp_functions_0_aMux_207_a2_combout;
wire fp_functions_0_aR_uid148_fpAddTest_q_a31_a_a0_combout;
wire fp_functions_0_arVStage_uid165_lzCountVal_uid85_fpAddTest_merged_bit_select_b_a2_a_a4_combout;
wire fp_functions_0_arVStage_uid165_lzCountVal_uid85_fpAddTest_merged_bit_select_b_a2_a_a5_combout;
wire fp_functions_0_arVStage_uid165_lzCountVal_uid85_fpAddTest_merged_bit_select_b_a3_a_a6_combout;
wire fp_functions_0_areduce_nor_6_a0_combout;
wire fp_functions_0_arVStage_uid165_lzCountVal_uid85_fpAddTest_merged_bit_select_b_a1_a_a7_combout;
wire fp_functions_0_areduce_nor_6_a1_combout;
wire fp_functions_0_arVStage_uid171_lzCountVal_uid85_fpAddTest_merged_bit_select_b_a1_a_a2_combout;
wire fp_functions_0_arVStage_uid171_lzCountVal_uid85_fpAddTest_merged_bit_select_b_a1_a_a3_combout;
wire fp_functions_0_arVStage_uid171_lzCountVal_uid85_fpAddTest_merged_bit_select_b_a0_a_a4_combout;
wire fp_functions_0_arVStage_uid171_lzCountVal_uid85_fpAddTest_merged_bit_select_b_a0_a_a5_combout;
wire fp_functions_0_areduce_nor_5_a0_combout;
wire fp_functions_0_arVStage_uid171_lzCountVal_uid85_fpAddTest_merged_bit_select_c_a1_a_a1_combout;
wire fp_functions_0_arVStage_uid171_lzCountVal_uid85_fpAddTest_merged_bit_select_c_a1_a_a2_combout;
wire fp_functions_0_arVStage_uid177_lzCountVal_uid85_fpAddTest_b_a0_a_a0_combout;
wire fp_functions_0_arVStage_uid177_lzCountVal_uid85_fpAddTest_b_a0_a_a1_combout;
wire fp_functions_0_areduce_nor_6_a2_combout;
wire fp_functions_0_areduce_nor_6_a3_combout;
wire fp_functions_0_areduce_nor_8_a0_combout;
wire fp_functions_0_areduce_nor_8_acombout;
wire fp_functions_0_areduce_nor_9_a0_combout;
wire fp_functions_0_areduce_nor_9_acombout;
wire fp_functions_0_aregInputs_uid118_fpAddTest_qi_a0_a_a1_combout;
wire fp_functions_0_aexcI_aSig_uid27_fpAddTest_q_a0_a_acombout;
wire fp_functions_0_aexcI_bSig_uid41_fpAddTest_q_a0_a_acombout;
wire fp_functions_0_aexcN_bSig_uid42_fpAddTest_qi_a0_a_acombout;
wire fp_functions_0_aexcN_aSig_uid28_fpAddTest_qi_a0_a_acombout;
wire fp_functions_0_asignRInfRZRReg_uid137_fpAddTest_qi_a0_a_a1_combout;
wire fp_functions_0_asignRInfRZRReg_uid137_fpAddTest_qi_a0_a_a2_combout;
wire fp_functions_0_ai2460_a1_combout;
wire fp_functions_0_ai2460_a2_combout;
wire fp_functions_0_ai2460_a3_combout;
wire fp_functions_0_areduce_nor_2_acombout;
wire fp_functions_0_ai2460_a4_combout;
wire fp_functions_0_ai2459_a1_combout;
wire fp_functions_0_ai2467_a0_combout;
wire fp_functions_0_ai2460_a5_combout;
wire fp_functions_0_ai2467_a1_combout;
wire fp_functions_0_ai2460_a6_combout;
wire fp_functions_0_ai2467_a2_combout;
wire fp_functions_0_ai2467_a3_combout;
wire fp_functions_0_ai2453_a1_combout;
wire fp_functions_0_ai2467_a4_combout;
wire fp_functions_0_ai2454_a1_combout;
wire fp_functions_0_ai2467_a5_combout;
wire fp_functions_0_ai2460_a7_combout;
wire fp_functions_0_ai2461_a1_combout;
wire fp_functions_0_ai2467_a6_combout;
wire fp_functions_0_ai2467_a7_combout;
wire fp_functions_0_ai2455_a1_combout;
wire fp_functions_0_ai2467_a8_combout;
wire fp_functions_0_ai2462_a1_combout;
wire fp_functions_0_ai2467_a9_combout;
wire fp_functions_0_ai2463_a1_combout;
wire fp_functions_0_ai2460_a8_combout;
wire fp_functions_0_ai2467_a10_combout;
wire fp_functions_0_areduce_nor_1_a0_combout;
wire fp_functions_0_areduce_nor_1_a1_combout;
wire fp_functions_0_areduce_nor_1_a2_combout;
wire fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a15_a_aq;
wire fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a14_a_aq;
wire fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a13_a_aq;
wire fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a12_a_aq;
wire fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a10_a_aq;
wire fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a11_a_aq;
wire fp_functions_0_areduce_nor_1_a3_combout;
wire fp_functions_0_areduce_nor_1_a4_combout;
wire fp_functions_0_ai2464_a1_combout;
wire fp_functions_0_ai2467_a11_combout;
wire fp_functions_0_ai2460_a9_combout;
wire fp_functions_0_ai2460_a10_combout;
wire fp_functions_0_ai2467_a12_combout;
wire fp_functions_0_ai2467_a13_combout;
wire fp_functions_0_ai2467_a14_combout;
wire fp_functions_0_ai2467_a15_combout;
wire fp_functions_0_afracBAddOpPostXor_uid81_fpAddTest_b_a26_a_acombout;
wire fp_functions_0_areduce_nor_11_a0_combout;
wire fp_functions_0_areduce_nor_11_a1_combout;
wire fp_functions_0_areduce_nor_11_a2_combout;
wire fp_functions_0_areduce_nor_11_a3_combout;
wire fp_functions_0_areduce_nor_11_a4_combout;
wire fp_functions_0_areduce_nor_11_acombout;
wire fp_functions_0_areduce_nor_4_acombout;
wire fp_functions_0_areduce_nor_3_acombout;
wire fp_functions_0_aMux_186_a0_combout;
wire fp_functions_0_aMux_186_a1_combout;
wire fp_functions_0_aMux_186_a2_combout;
wire fp_functions_0_ai3337_a0_combout;
wire fp_functions_0_areduce_nor_12_acombout;
wire fp_functions_0_aMux_186_a3_combout;
wire fp_functions_0_aMux_186_a4_combout;
wire fp_functions_0_ai3365_a0_combout;
wire fp_functions_0_aMux_186_a5_combout;
wire fp_functions_0_aMux_186_a6_combout;
wire fp_functions_0_ai3365_a1_combout;
wire fp_functions_0_aMux_186_a7_combout;
wire fp_functions_0_ai3365_a2_combout;
wire fp_functions_0_aMux_186_a8_combout;
wire fp_functions_0_aMux_186_a9_combout;
wire fp_functions_0_ai3365_a3_combout;
wire fp_functions_0_aMux_186_a10_combout;
wire fp_functions_0_aMux_186_a11_combout;
wire fp_functions_0_ai3365_a4_combout;
wire fp_functions_0_aMux_186_a12_combout;
wire fp_functions_0_aMux_186_a13_combout;
wire fp_functions_0_ai3365_a5_combout;
wire fp_functions_0_aMux_186_a14_combout;
wire fp_functions_0_aMux_186_a15_combout;
wire fp_functions_0_ai3365_a6_combout;
wire fp_functions_0_aMux_186_a16_combout;
wire fp_functions_0_aMux_186_a17_combout;
wire fp_functions_0_ai3365_a7_combout;
wire fp_functions_0_aMux_186_a18_combout;
wire fp_functions_0_aMux_186_a19_combout;
wire fp_functions_0_ai3365_a8_combout;
wire fp_functions_0_aMux_186_a20_combout;
wire fp_functions_0_aMux_186_a21_combout;
wire fp_functions_0_ai3365_a9_combout;
wire fp_functions_0_aMux_186_a22_combout;
wire fp_functions_0_aMux_186_a23_combout;
wire fp_functions_0_ai3365_a10_combout;
wire fp_functions_0_aMux_158_a0_combout;
wire fp_functions_0_aMux_186_a24_combout;
wire fp_functions_0_ai3365_a11_combout;
wire fp_functions_0_aMux_158_a1_combout;
wire fp_functions_0_aMux_186_a25_combout;
wire fp_functions_0_ai3365_a12_combout;
wire fp_functions_0_aMux_158_a2_combout;
wire fp_functions_0_aMux_186_a26_combout;
wire fp_functions_0_ai3365_a13_combout;
wire fp_functions_0_aMux_158_a3_combout;
wire fp_functions_0_aMux_186_a27_combout;
wire fp_functions_0_ai3365_a14_combout;
wire fp_functions_0_aMux_158_a4_combout;
wire fp_functions_0_aMux_186_a28_combout;
wire fp_functions_0_ai3365_a15_combout;
wire fp_functions_0_aMux_158_a5_combout;
wire fp_functions_0_aMux_186_a29_combout;
wire fp_functions_0_ai3365_a16_combout;
wire fp_functions_0_aMux_158_a6_combout;
wire fp_functions_0_aMux_186_a30_combout;
wire fp_functions_0_ai3365_a17_combout;
wire fp_functions_0_aMux_158_a7_combout;
wire fp_functions_0_aMux_186_a31_combout;
wire fp_functions_0_ai3337_a1_combout;
wire fp_functions_0_aMux_158_a8_combout;
wire fp_functions_0_aMux_186_a32_combout;
wire fp_functions_0_ai3365_a18_combout;
wire fp_functions_0_aMux_158_a9_combout;
wire fp_functions_0_aMux_186_a33_combout;
wire fp_functions_0_ai3365_a19_combout;
wire fp_functions_0_aMux_158_a10_combout;
wire fp_functions_0_aMux_186_a34_combout;
wire fp_functions_0_ai3337_a2_combout;
wire fp_functions_0_astickyBits_uid69_fpAddTest_merged_bit_select_b_a0_a_a0_combout;
wire fp_functions_0_astickyBits_uid69_fpAddTest_merged_bit_select_b_a0_a_a1_combout;
wire fp_functions_0_astickyBits_uid69_fpAddTest_merged_bit_select_b_a0_a_a2_combout;
wire fp_functions_0_astickyBits_uid69_fpAddTest_merged_bit_select_b_a0_a_a3_combout;
wire fp_functions_0_astickyBits_uid69_fpAddTest_merged_bit_select_b_a0_a_a4_combout;
wire fp_functions_0_astickyBits_uid69_fpAddTest_merged_bit_select_b_a0_a_a5_combout;
wire fp_functions_0_astickyBits_uid69_fpAddTest_merged_bit_select_b_a0_a_a6_combout;
wire fp_functions_0_astickyBits_uid69_fpAddTest_merged_bit_select_b_a0_a_a7_combout;
wire fp_functions_0_astickyBits_uid69_fpAddTest_merged_bit_select_b_a0_a_a8_combout;
wire fp_functions_0_astickyBits_uid69_fpAddTest_merged_bit_select_b_a0_a_a9_combout;
wire fp_functions_0_astickyBits_uid69_fpAddTest_merged_bit_select_b_a0_a_a10_combout;
wire fp_functions_0_astickyBits_uid69_fpAddTest_merged_bit_select_b_a0_a_a11_combout;
wire fp_functions_0_astickyBits_uid69_fpAddTest_merged_bit_select_b_a0_a_a12_combout;
wire fp_functions_0_astickyBits_uid69_fpAddTest_merged_bit_select_b_a0_a_a13_combout;
wire fp_functions_0_astickyBits_uid69_fpAddTest_merged_bit_select_b_a0_a_a14_combout;
wire fp_functions_0_astickyBits_uid69_fpAddTest_merged_bit_select_b_a0_a_a15_combout;
wire fp_functions_0_astickyBits_uid69_fpAddTest_merged_bit_select_b_a0_a_a16_combout;
wire fp_functions_0_astickyBits_uid69_fpAddTest_merged_bit_select_b_a0_a_a17_combout;
wire fp_functions_0_astickyBits_uid69_fpAddTest_merged_bit_select_b_a0_a_a18_combout;
wire fp_functions_0_astickyBits_uid69_fpAddTest_merged_bit_select_b_a0_a_a19_combout;
wire fp_functions_0_astickyBits_uid69_fpAddTest_merged_bit_select_b_a0_a_a20_combout;
wire fp_functions_0_astickyBits_uid69_fpAddTest_merged_bit_select_b_a0_a_a21_combout;
wire fp_functions_0_astickyBits_uid69_fpAddTest_merged_bit_select_b_a0_a_a22_combout;
wire fp_functions_0_astickyBits_uid69_fpAddTest_merged_bit_select_b_a0_a_a23_combout;
wire fp_functions_0_afrac_bSig_uid36_fpAddTest_b_a13_a_a0_combout;
wire fp_functions_0_afrac_bSig_uid36_fpAddTest_b_a14_a_a1_combout;
wire fp_functions_0_areduce_nor_0_a0_combout;
wire fp_functions_0_areduce_nor_0_a1_combout;
wire fp_functions_0_areduce_nor_0_a2_combout;
wire fp_functions_0_areduce_nor_0_a3_combout;
wire fp_functions_0_areduce_nor_0_acombout;
wire fp_functions_0_aMux_2_a0_combout;
wire fp_functions_0_afrac_bSig_uid36_fpAddTest_b_a15_a_a2_combout;
wire fp_functions_0_afrac_bSig_uid36_fpAddTest_b_a16_a_a3_combout;
wire fp_functions_0_aMux_2_a1_combout;
wire fp_functions_0_afrac_bSig_uid36_fpAddTest_b_a17_a_a4_combout;
wire fp_functions_0_afrac_bSig_uid36_fpAddTest_b_a18_a_a5_combout;
wire fp_functions_0_aMux_2_a2_combout;
wire fp_functions_0_afrac_bSig_uid36_fpAddTest_b_a19_a_a6_combout;
wire fp_functions_0_afrac_bSig_uid36_fpAddTest_b_a20_a_a7_combout;
wire fp_functions_0_aMux_2_a3_combout;
wire fp_functions_0_aMux_59_a0_combout;
wire fp_functions_0_afrac_bSig_uid36_fpAddTest_b_a5_a_a8_combout;
wire fp_functions_0_afrac_bSig_uid36_fpAddTest_b_a6_a_a9_combout;
wire fp_functions_0_aMux_2_a4_combout;
wire fp_functions_0_afrac_bSig_uid36_fpAddTest_b_a7_a_a10_combout;
wire fp_functions_0_afrac_bSig_uid36_fpAddTest_b_a8_a_a11_combout;
wire fp_functions_0_aMux_2_a5_combout;
wire fp_functions_0_afrac_bSig_uid36_fpAddTest_b_a9_a_a12_combout;
wire fp_functions_0_afrac_bSig_uid36_fpAddTest_b_a10_a_a13_combout;
wire fp_functions_0_aMux_2_a6_combout;
wire fp_functions_0_afrac_bSig_uid36_fpAddTest_b_a11_a_a14_combout;
wire fp_functions_0_afrac_bSig_uid36_fpAddTest_b_a12_a_a15_combout;
wire fp_functions_0_aMux_2_a7_combout;
wire fp_functions_0_aMux_59_a1_combout;
wire fp_functions_0_aMux_2_a8_combout;
wire fp_functions_0_aMux_2_a9_combout;
wire fp_functions_0_afrac_bSig_uid36_fpAddTest_b_a0_a_a16_combout;
wire fp_functions_0_aMux_2_a10_combout;
wire fp_functions_0_aMux_59_a2_combout;
wire fp_functions_0_afrac_bSig_uid36_fpAddTest_b_a21_a_a17_combout;
wire fp_functions_0_aMux_2_a11_combout;
wire fp_functions_0_afrac_bSig_uid36_fpAddTest_b_a22_a_a18_combout;
wire fp_functions_0_aMux_2_a12_combout;
wire fp_functions_0_aMux_59_a3_combout;
wire fp_functions_0_ai1783_a0_combout;
wire fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a28_a_a0_combout;
wire fp_functions_0_aMux_2_a13_combout;
wire fp_functions_0_aMux_57_a0_combout;
wire fp_functions_0_aMux_57_a1_combout;
wire fp_functions_0_aMux_65_a0_combout;
wire fp_functions_0_aMux_2_a14_combout;
wire fp_functions_0_aMux_2_a15_combout;
wire fp_functions_0_aMux_57_a2_combout;
wire fp_functions_0_aMux_49_a0_combout;
wire fp_functions_0_ai1734_a0_combout;
wire fp_functions_0_ai1734_a1_combout;
wire fp_functions_0_ai1734_a2_combout;
wire fp_functions_0_aMux_2_a16_combout;
wire fp_functions_0_aMux_2_a17_combout;
wire fp_functions_0_aMux_2_a18_combout;
wire fp_functions_0_aMux_2_a19_combout;
wire fp_functions_0_aMux_2_a20_combout;
wire fp_functions_0_aMux_60_a0_combout;
wire fp_functions_0_aMux_2_a21_combout;
wire fp_functions_0_aMux_2_a22_combout;
wire fp_functions_0_aMux_2_a23_combout;
wire fp_functions_0_aMux_2_a24_combout;
wire fp_functions_0_aMux_60_a1_combout;
wire fp_functions_0_aMux_23_a0_combout;
wire fp_functions_0_aMux_2_a25_combout;
wire fp_functions_0_aMux_2_a26_combout;
wire fp_functions_0_aMux_2_a27_combout;
wire fp_functions_0_aMux_23_a1_combout;
wire fp_functions_0_aMux_2_a28_combout;
wire fp_functions_0_aMux_2_a29_combout;
wire fp_functions_0_aMux_60_a2_combout;
wire fp_functions_0_ai1783_a1_combout;
wire fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a2_a_a1_combout;
wire fp_functions_0_ai1783_a2_combout;
wire fp_functions_0_aMux_57_a3_combout;
wire fp_functions_0_aMux_57_a4_combout;
wire fp_functions_0_aMux_61_a0_combout;
wire fp_functions_0_aMux_77_a0_combout;
wire fp_functions_0_ai1783_a3_combout;
wire fp_functions_0_aMux_60_a3_combout;
wire fp_functions_0_aMux_60_a4_combout;
wire fp_functions_0_aMux_76_a0_combout;
wire fp_functions_0_aMux_60_a5_combout;
wire fp_functions_0_ai1783_a4_combout;
wire fp_functions_0_ai1783_a5_combout;
wire fp_functions_0_aMux_58_a0_combout;
wire fp_functions_0_aMux_58_a1_combout;
wire fp_functions_0_aMux_78_a0_combout;
wire fp_functions_0_aMux_62_a0_combout;
wire fp_functions_0_ai1783_a6_combout;
wire fp_functions_0_ai1783_a7_combout;
wire fp_functions_0_aMux_59_a4_combout;
wire fp_functions_0_aMux_59_a5_combout;
wire fp_functions_0_aMux_59_a6_combout;
wire fp_functions_0_aMux_79_a0_combout;
wire fp_functions_0_ai1783_a8_combout;
wire fp_functions_0_aMux_57_a5_combout;
wire fp_functions_0_ai1783_a9_combout;
wire fp_functions_0_aMux_58_a2_combout;
wire fp_functions_0_aMux_58_a3_combout;
wire fp_functions_0_aMux_58_a4_combout;
wire fp_functions_0_ai1783_a10_combout;
wire fp_functions_0_ai1783_a11_combout;
wire fp_functions_0_ai1783_a12_combout;
wire fp_functions_0_ai1783_a13_combout;
wire fp_functions_0_ai1783_a14_combout;
wire fp_functions_0_ai1783_a15_combout;
wire fp_functions_0_aMux_50_a0_combout;
wire fp_functions_0_ai1783_a16_combout;
wire fp_functions_0_aMux_51_a0_combout;
wire fp_functions_0_ai1783_a17_combout;
wire fp_functions_0_aMux_52_a0_combout;
wire fp_functions_0_ai1783_a18_combout;
wire fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a13_a_a2_combout;
wire fp_functions_0_ai1783_a19_combout;
wire fp_functions_0_aMux_53_a1_combout;
wire fp_functions_0_aMux_54_a1_combout;
wire fp_functions_0_aexp_bSig_uid35_fpAddTest_b_a3_a_a0_combout;
wire fp_functions_0_aexp_bSig_uid35_fpAddTest_b_a1_a_a1_combout;
wire fp_functions_0_areduce_nor_7_a0_combout;
wire fp_functions_0_aexp_bSig_uid35_fpAddTest_b_a5_a_a2_combout;
wire fp_functions_0_areduce_nor_7_a1_combout;
wire fp_functions_0_aexp_bSig_uid35_fpAddTest_b_a7_a_a3_combout;
wire fp_functions_0_areduce_nor_7_a2_combout;
wire fp_functions_0_aexp_aSig_uid21_fpAddTest_b_a0_a_a0_combout;
wire fp_functions_0_aexp_aSig_uid21_fpAddTest_b_a0_a_a1_combout;
wire fp_functions_0_aexp_aSig_uid21_fpAddTest_b_a0_a_a2_combout;
wire fp_functions_0_aexp_aSig_uid21_fpAddTest_b_a0_a_a3_combout;
wire fp_functions_0_aexp_aSig_uid21_fpAddTest_b_a0_a_a4_combout;
wire fp_functions_0_aexp_aSig_uid21_fpAddTest_b_a0_a_a5_combout;
wire fp_functions_0_aexp_aSig_uid21_fpAddTest_b_a0_a_a6_combout;
wire fp_functions_0_aexp_aSig_uid21_fpAddTest_b_a0_a_a7_combout;
wire fp_functions_0_ai326_a0_combout;
wire fp_functions_0_ai289_a0_combout;
wire fp_functions_0_ai2131_a0_combout;
wire fp_functions_0_ai2131_a1_combout;
wire fp_functions_0_ai2131_a2_combout;
wire fp_functions_0_ai2131_a3_combout;
wire fp_functions_0_ai2131_a4_combout;
wire fp_functions_0_ai2131_a5_combout;
wire fp_functions_0_ai2131_a6_combout;
wire fp_functions_0_ai2131_a7_combout;
wire fp_functions_0_ai2131_a8_combout;
wire fp_functions_0_ai2131_a9_combout;
wire fp_functions_0_ai2131_a10_combout;
wire fp_functions_0_ai2131_a11_combout;
wire fp_functions_0_ai2131_a12_combout;
wire fp_functions_0_ai2131_a13_combout;
wire fp_functions_0_ai2131_a14_combout;
wire fp_functions_0_ai2131_a15_combout;
wire fp_functions_0_ai2131_a16_combout;
wire fp_functions_0_ai2131_a17_combout;
wire fp_functions_0_ai2131_a18_combout;
wire fp_functions_0_ai2131_a19_combout;
wire fp_functions_0_ai2131_a20_combout;
wire fp_functions_0_ai2131_a21_combout;
wire fp_functions_0_ai2131_a22_combout;
wire fp_functions_0_areduce_nor_10_a0_combout;
wire fp_functions_0_areduce_nor_10_a1_combout;
wire fp_functions_0_areduce_nor_10_a2_combout;
wire fp_functions_0_areduce_nor_10_a3_combout;
wire fp_functions_0_areduce_nor_10_a4_combout;
wire fp_functions_0_areduce_nor_10_a5_combout;
wire fp_functions_0_areduce_nor_10_a6_combout;
wire fp_functions_0_areduce_nor_10_a7_combout;
wire fp_functions_0_areduce_nor_10_a8_combout;
wire fp_functions_0_areduce_nor_10_acombout;
wire fp_functions_0_ai3337_a3_combout;
wire fp_functions_0_ai3337_a4_combout;
wire fp_functions_0_ai3337_a5_combout;
wire fp_functions_0_ai3337_a6_combout;
wire fp_functions_0_ai3337_a7_combout;
wire fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a41_a_a3_combout;
wire fp_functions_0_aMux_59_a7_combout;
wire fp_functions_0_aMux_63_a0_combout;
wire fp_functions_0_aMux_62_a1_combout;
wire fp_functions_0_aMux_61_a1_combout;
wire fp_functions_0_aMux_60_a6_combout;
wire fp_functions_0_aMux_58_a5_combout;
wire fp_functions_0_aMux_57_a6_combout;
wire fp_functions_0_aMux_56_a1_combout;
wire fp_functions_0_ai1783_a20_combout;
wire fp_functions_0_ai1783_a21_combout;
wire fp_functions_0_ai1783_a22_combout;
wire fp_functions_0_ai1783_a23_combout;
wire fp_functions_0_aMux_64_a0_combout;
wire fp_functions_0_ai1783_a24_combout;
wire fp_functions_0_ai1783_a25_combout;
wire fp_functions_0_ai1783_a26_combout;
wire fp_functions_0_ai1783_a27_combout;
wire fp_functions_0_ai1783_a28_combout;
wire fp_functions_0_ai1783_a29_combout;
wire fp_functions_0_ai1783_a30_combout;
wire fp_functions_0_ai1783_a31_combout;
wire fp_functions_0_ai1783_a32_combout;
wire fp_functions_0_ai1783_a33_combout;
wire fp_functions_0_areduce_nor_0_a_wirecell_combout;


fourteennm_ff fp_functions_0_aredist2_aMinusA_uid87_fpAddTest_q_1_q_a0_a(
	.clk(clk),
	.d(fp_functions_0_areduce_nor_6_a3_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist2_aMinusA_uid87_fpAddTest_q_1_q_a0_a_aq));
defparam fp_functions_0_aredist2_aMinusA_uid87_fpAddTest_q_1_q_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist2_aMinusA_uid87_fpAddTest_q_1_q_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aregInputs_uid118_fpAddTest_delay_adelay_signals_a0_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aregInputs_uid118_fpAddTest_qi_a0_a_a1_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aregInputs_uid118_fpAddTest_delay_adelay_signals_a0_a_a0_a_aq));
defparam fp_functions_0_aregInputs_uid118_fpAddTest_delay_adelay_signals_a0_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aregInputs_uid118_fpAddTest_delay_adelay_signals_a0_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist16_excZ_aSig_uid16_uid23_fpAddTest_q_1_q_a0_a(
	.clk(clk),
	.d(fp_functions_0_areduce_nor_9_acombout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist16_excZ_aSig_uid16_uid23_fpAddTest_q_1_q_a0_a_aq));
defparam fp_functions_0_aredist16_excZ_aSig_uid16_uid23_fpAddTest_q_1_q_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist16_excZ_aSig_uid16_uid23_fpAddTest_q_1_q_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist14_excZ_bSig_uid17_uid37_fpAddTest_q_3_q_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist13_excZ_bSig_uid17_uid37_fpAddTest_q_2_q_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist14_excZ_bSig_uid17_uid37_fpAddTest_q_3_q_a0_a_aq));
defparam fp_functions_0_aredist14_excZ_bSig_uid17_uid37_fpAddTest_q_3_q_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist14_excZ_bSig_uid17_uid37_fpAddTest_q_3_q_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist4_effSub_uid52_fpAddTest_q_2_q_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist4_effSub_uid52_fpAddTest_q_2_delay_0_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist4_effSub_uid52_fpAddTest_q_2_q_a0_a_aq));
defparam fp_functions_0_aredist4_effSub_uid52_fpAddTest_q_2_q_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist4_effSub_uid52_fpAddTest_q_2_q_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist15_excI_aSig_uid27_fpAddTest_q_1_q_a0_a(
	.clk(clk),
	.d(fp_functions_0_aexcI_aSig_uid27_fpAddTest_q_a0_a_acombout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist15_excI_aSig_uid27_fpAddTest_q_1_q_a0_a_aq));
defparam fp_functions_0_aredist15_excI_aSig_uid27_fpAddTest_q_1_q_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist15_excI_aSig_uid27_fpAddTest_q_1_q_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist10_excI_bSig_uid41_fpAddTest_q_1_q_a0_a(
	.clk(clk),
	.d(fp_functions_0_aexcI_bSig_uid41_fpAddTest_q_a0_a_acombout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist10_excI_bSig_uid41_fpAddTest_q_1_q_a0_a_aq));
defparam fp_functions_0_aredist10_excI_bSig_uid41_fpAddTest_q_1_q_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist10_excI_bSig_uid41_fpAddTest_q_1_q_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aexcN_bSig_uid42_fpAddTest_delay_adelay_signals_a0_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aexcN_bSig_uid42_fpAddTest_qi_a0_a_acombout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aexcN_bSig_uid42_fpAddTest_delay_adelay_signals_a0_a_a0_a_aq));
defparam fp_functions_0_aexcN_bSig_uid42_fpAddTest_delay_adelay_signals_a0_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aexcN_bSig_uid42_fpAddTest_delay_adelay_signals_a0_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aexcN_aSig_uid28_fpAddTest_delay_adelay_signals_a0_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_aexcN_aSig_uid28_fpAddTest_qi_a0_a_acombout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aexcN_aSig_uid28_fpAddTest_delay_adelay_signals_a0_a_a0_a_aq));
defparam fp_functions_0_aexcN_aSig_uid28_fpAddTest_delay_adelay_signals_a0_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aexcN_aSig_uid28_fpAddTest_delay_adelay_signals_a0_a_a0_a.power_up = "dont_care";

fourteennm_lcell_comb fp_functions_0_aadd_7_a1(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aleftShiftStage2_uid249_fracPostNormExt_uid88_fpAddTest_q_a4_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_7_a167_cout),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_7_a1_sumout),
	.cout(fp_functions_0_aadd_7_a2),
	.shareout());
defparam fp_functions_0_aadd_7_a1.extended_lut = "off";
defparam fp_functions_0_aadd_7_a1.lut_mask = 64'h0000000000000F0F;
defparam fp_functions_0_aadd_7_a1.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_7_a6(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aexpPostNorm_uid92_fpAddTest_o_a5_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_7_a32),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_7_a6_sumout),
	.cout(fp_functions_0_aadd_7_a7),
	.shareout());
defparam fp_functions_0_aadd_7_a6.extended_lut = "off";
defparam fp_functions_0_aadd_7_a6.lut_mask = 64'h0000000000000F0F;
defparam fp_functions_0_aadd_7_a6.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_7_a11(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aexpPostNorm_uid92_fpAddTest_o_a0_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_7_a162),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_7_a11_sumout),
	.cout(fp_functions_0_aadd_7_a12),
	.shareout());
defparam fp_functions_0_aadd_7_a11.extended_lut = "off";
defparam fp_functions_0_aadd_7_a11.lut_mask = 64'h0000000000000F0F;
defparam fp_functions_0_aadd_7_a11.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_7_a16(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aexpPostNorm_uid92_fpAddTest_o_a1_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_7_a12),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_7_a16_sumout),
	.cout(fp_functions_0_aadd_7_a17),
	.shareout());
defparam fp_functions_0_aadd_7_a16.extended_lut = "off";
defparam fp_functions_0_aadd_7_a16.lut_mask = 64'h0000000000000F0F;
defparam fp_functions_0_aadd_7_a16.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_7_a21(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aexpPostNorm_uid92_fpAddTest_o_a2_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_7_a17),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_7_a21_sumout),
	.cout(fp_functions_0_aadd_7_a22),
	.shareout());
defparam fp_functions_0_aadd_7_a21.extended_lut = "off";
defparam fp_functions_0_aadd_7_a21.lut_mask = 64'h0000000000000F0F;
defparam fp_functions_0_aadd_7_a21.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_7_a26(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aexpPostNorm_uid92_fpAddTest_o_a3_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_7_a22),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_7_a26_sumout),
	.cout(fp_functions_0_aadd_7_a27),
	.shareout());
defparam fp_functions_0_aadd_7_a26.extended_lut = "off";
defparam fp_functions_0_aadd_7_a26.lut_mask = 64'h0000000000000F0F;
defparam fp_functions_0_aadd_7_a26.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_7_a31(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aexpPostNorm_uid92_fpAddTest_o_a4_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_7_a27),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_7_a31_sumout),
	.cout(fp_functions_0_aadd_7_a32),
	.shareout());
defparam fp_functions_0_aadd_7_a31.extended_lut = "off";
defparam fp_functions_0_aadd_7_a31.lut_mask = 64'h0000000000000F0F;
defparam fp_functions_0_aadd_7_a31.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_7_a36(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aexpPostNorm_uid92_fpAddTest_o_a6_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_7_a7),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_7_a36_sumout),
	.cout(fp_functions_0_aadd_7_a37),
	.shareout());
defparam fp_functions_0_aadd_7_a36.extended_lut = "off";
defparam fp_functions_0_aadd_7_a36.lut_mask = 64'h0000000000000F0F;
defparam fp_functions_0_aadd_7_a36.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_7_a41(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aexpPostNorm_uid92_fpAddTest_o_a7_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_7_a37),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_7_a41_sumout),
	.cout(fp_functions_0_aadd_7_a42),
	.shareout());
defparam fp_functions_0_aadd_7_a41.extended_lut = "off";
defparam fp_functions_0_aadd_7_a41.lut_mask = 64'h0000000000000F0F;
defparam fp_functions_0_aadd_7_a41.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_7_a46(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aexpPostNorm_uid92_fpAddTest_o_a8_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_7_a42),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_7_a46_sumout),
	.cout(fp_functions_0_aadd_7_a47),
	.shareout());
defparam fp_functions_0_aadd_7_a46.extended_lut = "off";
defparam fp_functions_0_aadd_7_a46.lut_mask = 64'h0000000000000F0F;
defparam fp_functions_0_aadd_7_a46.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_7_a51(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aexpPostNorm_uid92_fpAddTest_o_a9_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_7_a47),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_7_a51_sumout),
	.cout(),
	.shareout());
defparam fp_functions_0_aadd_7_a51.extended_lut = "off";
defparam fp_functions_0_aadd_7_a51.lut_mask = 64'h0000000000000F0F;
defparam fp_functions_0_aadd_7_a51.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_7_a56(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aleftShiftStage2_uid249_fracPostNormExt_uid88_fpAddTest_q_a5_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_7_a2),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_7_a56_sumout),
	.cout(fp_functions_0_aadd_7_a57),
	.shareout());
defparam fp_functions_0_aadd_7_a56.extended_lut = "off";
defparam fp_functions_0_aadd_7_a56.lut_mask = 64'h0000000000000F0F;
defparam fp_functions_0_aadd_7_a56.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_7_a61(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aleftShiftStage2_uid249_fracPostNormExt_uid88_fpAddTest_q_a6_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_7_a57),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_7_a61_sumout),
	.cout(fp_functions_0_aadd_7_a62),
	.shareout());
defparam fp_functions_0_aadd_7_a61.extended_lut = "off";
defparam fp_functions_0_aadd_7_a61.lut_mask = 64'h0000000000000F0F;
defparam fp_functions_0_aadd_7_a61.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_7_a66(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aleftShiftStage2_uid249_fracPostNormExt_uid88_fpAddTest_q_a7_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_7_a62),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_7_a66_sumout),
	.cout(fp_functions_0_aadd_7_a67),
	.shareout());
defparam fp_functions_0_aadd_7_a66.extended_lut = "off";
defparam fp_functions_0_aadd_7_a66.lut_mask = 64'h0000000000000F0F;
defparam fp_functions_0_aadd_7_a66.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_7_a71(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aleftShiftStage2_uid249_fracPostNormExt_uid88_fpAddTest_q_a8_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_7_a67),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_7_a71_sumout),
	.cout(fp_functions_0_aadd_7_a72),
	.shareout());
defparam fp_functions_0_aadd_7_a71.extended_lut = "off";
defparam fp_functions_0_aadd_7_a71.lut_mask = 64'h0000000000000F0F;
defparam fp_functions_0_aadd_7_a71.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_7_a76(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aleftShiftStage2_uid249_fracPostNormExt_uid88_fpAddTest_q_a9_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_7_a72),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_7_a76_sumout),
	.cout(fp_functions_0_aadd_7_a77),
	.shareout());
defparam fp_functions_0_aadd_7_a76.extended_lut = "off";
defparam fp_functions_0_aadd_7_a76.lut_mask = 64'h0000000000000F0F;
defparam fp_functions_0_aadd_7_a76.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_7_a81(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aleftShiftStage2_uid249_fracPostNormExt_uid88_fpAddTest_q_a10_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_7_a77),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_7_a81_sumout),
	.cout(fp_functions_0_aadd_7_a82),
	.shareout());
defparam fp_functions_0_aadd_7_a81.extended_lut = "off";
defparam fp_functions_0_aadd_7_a81.lut_mask = 64'h0000000000000F0F;
defparam fp_functions_0_aadd_7_a81.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_7_a86(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aleftShiftStage2_uid249_fracPostNormExt_uid88_fpAddTest_q_a11_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_7_a82),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_7_a86_sumout),
	.cout(fp_functions_0_aadd_7_a87),
	.shareout());
defparam fp_functions_0_aadd_7_a86.extended_lut = "off";
defparam fp_functions_0_aadd_7_a86.lut_mask = 64'h0000000000000F0F;
defparam fp_functions_0_aadd_7_a86.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_7_a91(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aleftShiftStage2_uid249_fracPostNormExt_uid88_fpAddTest_q_a12_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_7_a87),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_7_a91_sumout),
	.cout(fp_functions_0_aadd_7_a92),
	.shareout());
defparam fp_functions_0_aadd_7_a91.extended_lut = "off";
defparam fp_functions_0_aadd_7_a91.lut_mask = 64'h0000000000000F0F;
defparam fp_functions_0_aadd_7_a91.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_7_a96(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aleftShiftStage2_uid249_fracPostNormExt_uid88_fpAddTest_q_a13_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_7_a92),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_7_a96_sumout),
	.cout(fp_functions_0_aadd_7_a97),
	.shareout());
defparam fp_functions_0_aadd_7_a96.extended_lut = "off";
defparam fp_functions_0_aadd_7_a96.lut_mask = 64'h0000000000000F0F;
defparam fp_functions_0_aadd_7_a96.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_7_a101(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aleftShiftStage2_uid249_fracPostNormExt_uid88_fpAddTest_q_a14_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_7_a97),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_7_a101_sumout),
	.cout(fp_functions_0_aadd_7_a102),
	.shareout());
defparam fp_functions_0_aadd_7_a101.extended_lut = "off";
defparam fp_functions_0_aadd_7_a101.lut_mask = 64'h0000000000000F0F;
defparam fp_functions_0_aadd_7_a101.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_7_a106(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aleftShiftStage2_uid249_fracPostNormExt_uid88_fpAddTest_q_a15_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_7_a102),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_7_a106_sumout),
	.cout(fp_functions_0_aadd_7_a107),
	.shareout());
defparam fp_functions_0_aadd_7_a106.extended_lut = "off";
defparam fp_functions_0_aadd_7_a106.lut_mask = 64'h0000000000000F0F;
defparam fp_functions_0_aadd_7_a106.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_7_a111(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aleftShiftStage2_uid249_fracPostNormExt_uid88_fpAddTest_q_a16_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_7_a107),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_7_a111_sumout),
	.cout(fp_functions_0_aadd_7_a112),
	.shareout());
defparam fp_functions_0_aadd_7_a111.extended_lut = "off";
defparam fp_functions_0_aadd_7_a111.lut_mask = 64'h0000000000000F0F;
defparam fp_functions_0_aadd_7_a111.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_7_a116(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aleftShiftStage2_uid249_fracPostNormExt_uid88_fpAddTest_q_a17_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_7_a112),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_7_a116_sumout),
	.cout(fp_functions_0_aadd_7_a117),
	.shareout());
defparam fp_functions_0_aadd_7_a116.extended_lut = "off";
defparam fp_functions_0_aadd_7_a116.lut_mask = 64'h0000000000000F0F;
defparam fp_functions_0_aadd_7_a116.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_7_a121(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aleftShiftStage2_uid249_fracPostNormExt_uid88_fpAddTest_q_a18_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_7_a117),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_7_a121_sumout),
	.cout(fp_functions_0_aadd_7_a122),
	.shareout());
defparam fp_functions_0_aadd_7_a121.extended_lut = "off";
defparam fp_functions_0_aadd_7_a121.lut_mask = 64'h0000000000000F0F;
defparam fp_functions_0_aadd_7_a121.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_7_a126(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aleftShiftStage2_uid249_fracPostNormExt_uid88_fpAddTest_q_a19_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_7_a122),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_7_a126_sumout),
	.cout(fp_functions_0_aadd_7_a127),
	.shareout());
defparam fp_functions_0_aadd_7_a126.extended_lut = "off";
defparam fp_functions_0_aadd_7_a126.lut_mask = 64'h0000000000000F0F;
defparam fp_functions_0_aadd_7_a126.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_7_a131(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aleftShiftStage2_uid249_fracPostNormExt_uid88_fpAddTest_q_a20_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_7_a127),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_7_a131_sumout),
	.cout(fp_functions_0_aadd_7_a132),
	.shareout());
defparam fp_functions_0_aadd_7_a131.extended_lut = "off";
defparam fp_functions_0_aadd_7_a131.lut_mask = 64'h0000000000000F0F;
defparam fp_functions_0_aadd_7_a131.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_7_a136(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aleftShiftStage2_uid249_fracPostNormExt_uid88_fpAddTest_q_a21_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_7_a132),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_7_a136_sumout),
	.cout(fp_functions_0_aadd_7_a137),
	.shareout());
defparam fp_functions_0_aadd_7_a136.extended_lut = "off";
defparam fp_functions_0_aadd_7_a136.lut_mask = 64'h0000000000000F0F;
defparam fp_functions_0_aadd_7_a136.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_7_a141(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aleftShiftStage2_uid249_fracPostNormExt_uid88_fpAddTest_q_a22_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_7_a137),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_7_a141_sumout),
	.cout(fp_functions_0_aadd_7_a142),
	.shareout());
defparam fp_functions_0_aadd_7_a141.extended_lut = "off";
defparam fp_functions_0_aadd_7_a141.lut_mask = 64'h0000000000000F0F;
defparam fp_functions_0_aadd_7_a141.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_7_a146(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aleftShiftStage2_uid249_fracPostNormExt_uid88_fpAddTest_q_a23_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_7_a142),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_7_a146_sumout),
	.cout(fp_functions_0_aadd_7_a147),
	.shareout());
defparam fp_functions_0_aadd_7_a146.extended_lut = "off";
defparam fp_functions_0_aadd_7_a146.lut_mask = 64'h0000000000000F0F;
defparam fp_functions_0_aadd_7_a146.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_7_a151(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aleftShiftStage2_uid249_fracPostNormExt_uid88_fpAddTest_q_a24_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_7_a147),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_7_a151_sumout),
	.cout(fp_functions_0_aadd_7_a152),
	.shareout());
defparam fp_functions_0_aadd_7_a151.extended_lut = "off";
defparam fp_functions_0_aadd_7_a151.lut_mask = 64'h0000000000000F0F;
defparam fp_functions_0_aadd_7_a151.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_7_a156(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aleftShiftStage2_uid249_fracPostNormExt_uid88_fpAddTest_q_a25_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_7_a152),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_7_a156_sumout),
	.cout(fp_functions_0_aadd_7_a157),
	.shareout());
defparam fp_functions_0_aadd_7_a156.extended_lut = "off";
defparam fp_functions_0_aadd_7_a156.lut_mask = 64'h0000000000000F0F;
defparam fp_functions_0_aadd_7_a156.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_7_a161(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aleftShiftStage2_uid249_fracPostNormExt_uid88_fpAddTest_q_a26_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_7_a157),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_7_a161_sumout),
	.cout(fp_functions_0_aadd_7_a162),
	.shareout());
defparam fp_functions_0_aadd_7_a161.extended_lut = "off";
defparam fp_functions_0_aadd_7_a161.lut_mask = 64'h0000000000000F0F;
defparam fp_functions_0_aadd_7_a161.shared_arith = "off";

fourteennm_ff fp_functions_0_asignRInfRZRReg_uid137_fpAddTest_delay_adelay_signals_a0_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_asignRInfRZRReg_uid137_fpAddTest_qi_a0_a_a2_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_asignRInfRZRReg_uid137_fpAddTest_delay_adelay_signals_a0_a_a0_a_aq));
defparam fp_functions_0_asignRInfRZRReg_uid137_fpAddTest_delay_adelay_signals_a0_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_asignRInfRZRReg_uid137_fpAddTest_delay_adelay_signals_a0_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist1_vCount_uid152_lzCountVal_uid85_fpAddTest_q_1_q_a0_a(
	.clk(clk),
	.d(fp_functions_0_areduce_nor_2_acombout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist1_vCount_uid152_lzCountVal_uid85_fpAddTest_q_1_q_a0_a_aq));
defparam fp_functions_0_aredist1_vCount_uid152_lzCountVal_uid85_fpAddTest_q_1_q_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist1_vCount_uid152_lzCountVal_uid85_fpAddTest_q_1_q_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_avStagei_uid157_lzCountVal_uid85_fpAddTest_q_a11_a(
	.clk(clk),
	.d(fp_functions_0_ai2467_a0_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_avStagei_uid157_lzCountVal_uid85_fpAddTest_q_a11_a_aq));
defparam fp_functions_0_avStagei_uid157_lzCountVal_uid85_fpAddTest_q_a11_a.is_wysiwyg = "true";
defparam fp_functions_0_avStagei_uid157_lzCountVal_uid85_fpAddTest_q_a11_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_avStagei_uid157_lzCountVal_uid85_fpAddTest_q_a10_a(
	.clk(clk),
	.d(fp_functions_0_ai2467_a1_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_avStagei_uid157_lzCountVal_uid85_fpAddTest_q_a10_a_aq));
defparam fp_functions_0_avStagei_uid157_lzCountVal_uid85_fpAddTest_q_a10_a.is_wysiwyg = "true";
defparam fp_functions_0_avStagei_uid157_lzCountVal_uid85_fpAddTest_q_a10_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_avStagei_uid157_lzCountVal_uid85_fpAddTest_q_a8_a(
	.clk(clk),
	.d(fp_functions_0_ai2467_a2_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_avStagei_uid157_lzCountVal_uid85_fpAddTest_q_a8_a_aq));
defparam fp_functions_0_avStagei_uid157_lzCountVal_uid85_fpAddTest_q_a8_a.is_wysiwyg = "true";
defparam fp_functions_0_avStagei_uid157_lzCountVal_uid85_fpAddTest_q_a8_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_avStagei_uid157_lzCountVal_uid85_fpAddTest_q_a9_a(
	.clk(clk),
	.d(fp_functions_0_ai2467_a3_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_avStagei_uid157_lzCountVal_uid85_fpAddTest_q_a9_a_aq));
defparam fp_functions_0_avStagei_uid157_lzCountVal_uid85_fpAddTest_q_a9_a.is_wysiwyg = "true";
defparam fp_functions_0_avStagei_uid157_lzCountVal_uid85_fpAddTest_q_a9_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_avStagei_uid157_lzCountVal_uid85_fpAddTest_q_a15_a(
	.clk(clk),
	.d(fp_functions_0_ai2467_a4_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_avStagei_uid157_lzCountVal_uid85_fpAddTest_q_a15_a_aq));
defparam fp_functions_0_avStagei_uid157_lzCountVal_uid85_fpAddTest_q_a15_a.is_wysiwyg = "true";
defparam fp_functions_0_avStagei_uid157_lzCountVal_uid85_fpAddTest_q_a15_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_avStagei_uid157_lzCountVal_uid85_fpAddTest_q_a14_a(
	.clk(clk),
	.d(fp_functions_0_ai2467_a5_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_avStagei_uid157_lzCountVal_uid85_fpAddTest_q_a14_a_aq));
defparam fp_functions_0_avStagei_uid157_lzCountVal_uid85_fpAddTest_q_a14_a.is_wysiwyg = "true";
defparam fp_functions_0_avStagei_uid157_lzCountVal_uid85_fpAddTest_q_a14_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_avStagei_uid157_lzCountVal_uid85_fpAddTest_q_a7_a(
	.clk(clk),
	.d(fp_functions_0_ai2467_a6_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_avStagei_uid157_lzCountVal_uid85_fpAddTest_q_a7_a_aq));
defparam fp_functions_0_avStagei_uid157_lzCountVal_uid85_fpAddTest_q_a7_a.is_wysiwyg = "true";
defparam fp_functions_0_avStagei_uid157_lzCountVal_uid85_fpAddTest_q_a7_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_avStagei_uid157_lzCountVal_uid85_fpAddTest_q_a12_a(
	.clk(clk),
	.d(fp_functions_0_ai2467_a7_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_avStagei_uid157_lzCountVal_uid85_fpAddTest_q_a12_a_aq));
defparam fp_functions_0_avStagei_uid157_lzCountVal_uid85_fpAddTest_q_a12_a.is_wysiwyg = "true";
defparam fp_functions_0_avStagei_uid157_lzCountVal_uid85_fpAddTest_q_a12_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_avStagei_uid157_lzCountVal_uid85_fpAddTest_q_a13_a(
	.clk(clk),
	.d(fp_functions_0_ai2467_a8_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_avStagei_uid157_lzCountVal_uid85_fpAddTest_q_a13_a_aq));
defparam fp_functions_0_avStagei_uid157_lzCountVal_uid85_fpAddTest_q_a13_a.is_wysiwyg = "true";
defparam fp_functions_0_avStagei_uid157_lzCountVal_uid85_fpAddTest_q_a13_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_avStagei_uid157_lzCountVal_uid85_fpAddTest_q_a6_a(
	.clk(clk),
	.d(fp_functions_0_ai2467_a9_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_avStagei_uid157_lzCountVal_uid85_fpAddTest_q_a6_a_aq));
defparam fp_functions_0_avStagei_uid157_lzCountVal_uid85_fpAddTest_q_a6_a.is_wysiwyg = "true";
defparam fp_functions_0_avStagei_uid157_lzCountVal_uid85_fpAddTest_q_a6_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_avStagei_uid157_lzCountVal_uid85_fpAddTest_q_a5_a(
	.clk(clk),
	.d(fp_functions_0_ai2467_a10_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_avStagei_uid157_lzCountVal_uid85_fpAddTest_q_a5_a_aq));
defparam fp_functions_0_avStagei_uid157_lzCountVal_uid85_fpAddTest_q_a5_a.is_wysiwyg = "true";
defparam fp_functions_0_avStagei_uid157_lzCountVal_uid85_fpAddTest_q_a5_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_avStagei_uid157_lzCountVal_uid85_fpAddTest_q_a4_a(
	.clk(clk),
	.d(fp_functions_0_ai2467_a11_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_avStagei_uid157_lzCountVal_uid85_fpAddTest_q_a4_a_aq));
defparam fp_functions_0_avStagei_uid157_lzCountVal_uid85_fpAddTest_q_a4_a.is_wysiwyg = "true";
defparam fp_functions_0_avStagei_uid157_lzCountVal_uid85_fpAddTest_q_a4_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_avStagei_uid157_lzCountVal_uid85_fpAddTest_q_a3_a(
	.clk(clk),
	.d(fp_functions_0_ai2467_a12_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_avStagei_uid157_lzCountVal_uid85_fpAddTest_q_a3_a_aq));
defparam fp_functions_0_avStagei_uid157_lzCountVal_uid85_fpAddTest_q_a3_a.is_wysiwyg = "true";
defparam fp_functions_0_avStagei_uid157_lzCountVal_uid85_fpAddTest_q_a3_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_avStagei_uid157_lzCountVal_uid85_fpAddTest_q_a2_a(
	.clk(clk),
	.d(fp_functions_0_ai2467_a13_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_avStagei_uid157_lzCountVal_uid85_fpAddTest_q_a2_a_aq));
defparam fp_functions_0_avStagei_uid157_lzCountVal_uid85_fpAddTest_q_a2_a.is_wysiwyg = "true";
defparam fp_functions_0_avStagei_uid157_lzCountVal_uid85_fpAddTest_q_a2_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_avStagei_uid157_lzCountVal_uid85_fpAddTest_q_a1_a(
	.clk(clk),
	.d(fp_functions_0_ai2467_a15_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_avStagei_uid157_lzCountVal_uid85_fpAddTest_q_a1_a_aq));
defparam fp_functions_0_avStagei_uid157_lzCountVal_uid85_fpAddTest_q_a1_a.is_wysiwyg = "true";
defparam fp_functions_0_avStagei_uid157_lzCountVal_uid85_fpAddTest_q_a1_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist12_expXIsMax_uid38_fpAddTest_q_2_q_a0_a(
	.clk(clk),
	.d(fp_functions_0_aexpXIsMax_uid38_fpAddTest_delay_adelay_signals_a0_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist12_expXIsMax_uid38_fpAddTest_q_2_q_a0_a_aq));
defparam fp_functions_0_aredist12_expXIsMax_uid38_fpAddTest_q_2_q_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist12_expXIsMax_uid38_fpAddTest_q_2_q_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist9_InvExpXIsZero_uid44_fpAddTest_q_2_q_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist9_InvExpXIsZero_uid44_fpAddTest_q_2_delay_0_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist9_InvExpXIsZero_uid44_fpAddTest_q_2_q_a0_a_aq));
defparam fp_functions_0_aredist9_InvExpXIsZero_uid44_fpAddTest_q_2_q_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist9_InvExpXIsZero_uid44_fpAddTest_q_2_q_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist18_exp_aSig_uid21_fpAddTest_b_2_q_a4_a(
	.clk(clk),
	.d(fp_functions_0_aredist18_exp_aSig_uid21_fpAddTest_b_2_delay_0_a4_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist18_exp_aSig_uid21_fpAddTest_b_2_q_a4_a_aq));
defparam fp_functions_0_aredist18_exp_aSig_uid21_fpAddTest_b_2_q_a4_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist18_exp_aSig_uid21_fpAddTest_b_2_q_a4_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist18_exp_aSig_uid21_fpAddTest_b_2_q_a5_a(
	.clk(clk),
	.d(fp_functions_0_aredist18_exp_aSig_uid21_fpAddTest_b_2_delay_0_a5_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist18_exp_aSig_uid21_fpAddTest_b_2_q_a5_a_aq));
defparam fp_functions_0_aredist18_exp_aSig_uid21_fpAddTest_b_2_q_a5_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist18_exp_aSig_uid21_fpAddTest_b_2_q_a5_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist18_exp_aSig_uid21_fpAddTest_b_2_q_a6_a(
	.clk(clk),
	.d(fp_functions_0_aredist18_exp_aSig_uid21_fpAddTest_b_2_delay_0_a6_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist18_exp_aSig_uid21_fpAddTest_b_2_q_a6_a_aq));
defparam fp_functions_0_aredist18_exp_aSig_uid21_fpAddTest_b_2_q_a6_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist18_exp_aSig_uid21_fpAddTest_b_2_q_a6_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist18_exp_aSig_uid21_fpAddTest_b_2_q_a7_a(
	.clk(clk),
	.d(fp_functions_0_aredist18_exp_aSig_uid21_fpAddTest_b_2_delay_0_a7_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist18_exp_aSig_uid21_fpAddTest_b_2_q_a7_a_aq));
defparam fp_functions_0_aredist18_exp_aSig_uid21_fpAddTest_b_2_q_a7_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist18_exp_aSig_uid21_fpAddTest_b_2_q_a7_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist18_exp_aSig_uid21_fpAddTest_b_2_q_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist18_exp_aSig_uid21_fpAddTest_b_2_delay_0_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist18_exp_aSig_uid21_fpAddTest_b_2_q_a0_a_aq));
defparam fp_functions_0_aredist18_exp_aSig_uid21_fpAddTest_b_2_q_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist18_exp_aSig_uid21_fpAddTest_b_2_q_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist18_exp_aSig_uid21_fpAddTest_b_2_q_a1_a(
	.clk(clk),
	.d(fp_functions_0_aredist18_exp_aSig_uid21_fpAddTest_b_2_delay_0_a1_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist18_exp_aSig_uid21_fpAddTest_b_2_q_a1_a_aq));
defparam fp_functions_0_aredist18_exp_aSig_uid21_fpAddTest_b_2_q_a1_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist18_exp_aSig_uid21_fpAddTest_b_2_q_a1_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist18_exp_aSig_uid21_fpAddTest_b_2_q_a2_a(
	.clk(clk),
	.d(fp_functions_0_aredist18_exp_aSig_uid21_fpAddTest_b_2_delay_0_a2_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist18_exp_aSig_uid21_fpAddTest_b_2_q_a2_a_aq));
defparam fp_functions_0_aredist18_exp_aSig_uid21_fpAddTest_b_2_q_a2_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist18_exp_aSig_uid21_fpAddTest_b_2_q_a2_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist18_exp_aSig_uid21_fpAddTest_b_2_q_a3_a(
	.clk(clk),
	.d(fp_functions_0_aredist18_exp_aSig_uid21_fpAddTest_b_2_delay_0_a3_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist18_exp_aSig_uid21_fpAddTest_b_2_q_a3_a_aq));
defparam fp_functions_0_aredist18_exp_aSig_uid21_fpAddTest_b_2_q_a3_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist18_exp_aSig_uid21_fpAddTest_b_2_q_a3_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist13_excZ_bSig_uid17_uid37_fpAddTest_q_2_q_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist13_excZ_bSig_uid17_uid37_fpAddTest_q_2_delay_0_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist13_excZ_bSig_uid17_uid37_fpAddTest_q_2_q_a0_a_aq));
defparam fp_functions_0_aredist13_excZ_bSig_uid17_uid37_fpAddTest_q_2_q_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist13_excZ_bSig_uid17_uid37_fpAddTest_q_2_q_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist4_effSub_uid52_fpAddTest_q_2_delay_0_a0_a(
	.clk(clk),
	.d(fp_functions_0_afracBAddOpPostXor_uid81_fpAddTest_b_a26_a_acombout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist4_effSub_uid52_fpAddTest_q_2_delay_0_a0_a_aq));
defparam fp_functions_0_aredist4_effSub_uid52_fpAddTest_q_2_delay_0_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist4_effSub_uid52_fpAddTest_q_2_delay_0_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_afracXIsZero_uid25_fpAddTest_delay_adelay_signals_a0_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_areduce_nor_11_acombout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_afracXIsZero_uid25_fpAddTest_delay_adelay_signals_a0_a_a0_a_aq));
defparam fp_functions_0_afracXIsZero_uid25_fpAddTest_delay_adelay_signals_a0_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_afracXIsZero_uid25_fpAddTest_delay_adelay_signals_a0_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist11_fracXIsZero_uid39_fpAddTest_q_2_q_a0_a(
	.clk(clk),
	.d(fp_functions_0_afracXIsZero_uid39_fpAddTest_delay_adelay_signals_a0_a_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist11_fracXIsZero_uid39_fpAddTest_q_2_q_a0_a_aq));
defparam fp_functions_0_aredist11_fracXIsZero_uid39_fpAddTest_q_2_q_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist11_fracXIsZero_uid39_fpAddTest_q_2_q_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aleftShiftStage2_uid249_fracPostNormExt_uid88_fpAddTest_q_a4_a(
	.clk(clk),
	.d(fp_functions_0_ai3337_a0_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aleftShiftStage2_uid249_fracPostNormExt_uid88_fpAddTest_q_a4_a_aq));
defparam fp_functions_0_aleftShiftStage2_uid249_fracPostNormExt_uid88_fpAddTest_q_a4_a.is_wysiwyg = "true";
defparam fp_functions_0_aleftShiftStage2_uid249_fracPostNormExt_uid88_fpAddTest_q_a4_a.power_up = "dont_care";

fourteennm_lcell_comb fp_functions_0_aadd_7_a167(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aleftShiftStage2_uid249_fracPostNormExt_uid88_fpAddTest_q_a3_a_aq),
	.datad(!fp_functions_0_areduce_nor_12_acombout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fp_functions_0_aadd_7_a167_cout),
	.shareout());
defparam fp_functions_0_aadd_7_a167.extended_lut = "off";
defparam fp_functions_0_aadd_7_a167.lut_mask = 64'h00000000000F0FF0;
defparam fp_functions_0_aadd_7_a167.shared_arith = "off";

fourteennm_ff fp_functions_0_aexpPostNorm_uid92_fpAddTest_o_a5_a(
	.clk(clk),
	.d(fp_functions_0_aadd_6_a1_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aexpPostNorm_uid92_fpAddTest_o_a5_a_aq));
defparam fp_functions_0_aexpPostNorm_uid92_fpAddTest_o_a5_a.is_wysiwyg = "true";
defparam fp_functions_0_aexpPostNorm_uid92_fpAddTest_o_a5_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aexpPostNorm_uid92_fpAddTest_o_a0_a(
	.clk(clk),
	.d(fp_functions_0_aadd_6_a6_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aexpPostNorm_uid92_fpAddTest_o_a0_a_aq));
defparam fp_functions_0_aexpPostNorm_uid92_fpAddTest_o_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aexpPostNorm_uid92_fpAddTest_o_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aexpPostNorm_uid92_fpAddTest_o_a1_a(
	.clk(clk),
	.d(fp_functions_0_aadd_6_a11_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aexpPostNorm_uid92_fpAddTest_o_a1_a_aq));
defparam fp_functions_0_aexpPostNorm_uid92_fpAddTest_o_a1_a.is_wysiwyg = "true";
defparam fp_functions_0_aexpPostNorm_uid92_fpAddTest_o_a1_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aexpPostNorm_uid92_fpAddTest_o_a2_a(
	.clk(clk),
	.d(fp_functions_0_aadd_6_a16_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aexpPostNorm_uid92_fpAddTest_o_a2_a_aq));
defparam fp_functions_0_aexpPostNorm_uid92_fpAddTest_o_a2_a.is_wysiwyg = "true";
defparam fp_functions_0_aexpPostNorm_uid92_fpAddTest_o_a2_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aexpPostNorm_uid92_fpAddTest_o_a3_a(
	.clk(clk),
	.d(fp_functions_0_aadd_6_a21_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aexpPostNorm_uid92_fpAddTest_o_a3_a_aq));
defparam fp_functions_0_aexpPostNorm_uid92_fpAddTest_o_a3_a.is_wysiwyg = "true";
defparam fp_functions_0_aexpPostNorm_uid92_fpAddTest_o_a3_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aexpPostNorm_uid92_fpAddTest_o_a4_a(
	.clk(clk),
	.d(fp_functions_0_aadd_6_a26_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aexpPostNorm_uid92_fpAddTest_o_a4_a_aq));
defparam fp_functions_0_aexpPostNorm_uid92_fpAddTest_o_a4_a.is_wysiwyg = "true";
defparam fp_functions_0_aexpPostNorm_uid92_fpAddTest_o_a4_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aexpPostNorm_uid92_fpAddTest_o_a6_a(
	.clk(clk),
	.d(fp_functions_0_aadd_6_a31_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aexpPostNorm_uid92_fpAddTest_o_a6_a_aq));
defparam fp_functions_0_aexpPostNorm_uid92_fpAddTest_o_a6_a.is_wysiwyg = "true";
defparam fp_functions_0_aexpPostNorm_uid92_fpAddTest_o_a6_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aexpPostNorm_uid92_fpAddTest_o_a7_a(
	.clk(clk),
	.d(fp_functions_0_aadd_6_a36_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aexpPostNorm_uid92_fpAddTest_o_a7_a_aq));
defparam fp_functions_0_aexpPostNorm_uid92_fpAddTest_o_a7_a.is_wysiwyg = "true";
defparam fp_functions_0_aexpPostNorm_uid92_fpAddTest_o_a7_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aexpPostNorm_uid92_fpAddTest_o_a8_a(
	.clk(clk),
	.d(fp_functions_0_aadd_6_a41_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aexpPostNorm_uid92_fpAddTest_o_a8_a_aq));
defparam fp_functions_0_aexpPostNorm_uid92_fpAddTest_o_a8_a.is_wysiwyg = "true";
defparam fp_functions_0_aexpPostNorm_uid92_fpAddTest_o_a8_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aexpPostNorm_uid92_fpAddTest_o_a9_a(
	.clk(clk),
	.d(fp_functions_0_aadd_6_a46_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aexpPostNorm_uid92_fpAddTest_o_a9_a_aq));
defparam fp_functions_0_aexpPostNorm_uid92_fpAddTest_o_a9_a.is_wysiwyg = "true";
defparam fp_functions_0_aexpPostNorm_uid92_fpAddTest_o_a9_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aleftShiftStage2_uid249_fracPostNormExt_uid88_fpAddTest_q_a5_a(
	.clk(clk),
	.d(fp_functions_0_ai3365_a0_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aleftShiftStage2_uid249_fracPostNormExt_uid88_fpAddTest_q_a5_a_aq));
defparam fp_functions_0_aleftShiftStage2_uid249_fracPostNormExt_uid88_fpAddTest_q_a5_a.is_wysiwyg = "true";
defparam fp_functions_0_aleftShiftStage2_uid249_fracPostNormExt_uid88_fpAddTest_q_a5_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aleftShiftStage2_uid249_fracPostNormExt_uid88_fpAddTest_q_a6_a(
	.clk(clk),
	.d(fp_functions_0_ai3365_a1_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aleftShiftStage2_uid249_fracPostNormExt_uid88_fpAddTest_q_a6_a_aq));
defparam fp_functions_0_aleftShiftStage2_uid249_fracPostNormExt_uid88_fpAddTest_q_a6_a.is_wysiwyg = "true";
defparam fp_functions_0_aleftShiftStage2_uid249_fracPostNormExt_uid88_fpAddTest_q_a6_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aleftShiftStage2_uid249_fracPostNormExt_uid88_fpAddTest_q_a7_a(
	.clk(clk),
	.d(fp_functions_0_ai3365_a2_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aleftShiftStage2_uid249_fracPostNormExt_uid88_fpAddTest_q_a7_a_aq));
defparam fp_functions_0_aleftShiftStage2_uid249_fracPostNormExt_uid88_fpAddTest_q_a7_a.is_wysiwyg = "true";
defparam fp_functions_0_aleftShiftStage2_uid249_fracPostNormExt_uid88_fpAddTest_q_a7_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aleftShiftStage2_uid249_fracPostNormExt_uid88_fpAddTest_q_a8_a(
	.clk(clk),
	.d(fp_functions_0_ai3365_a3_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aleftShiftStage2_uid249_fracPostNormExt_uid88_fpAddTest_q_a8_a_aq));
defparam fp_functions_0_aleftShiftStage2_uid249_fracPostNormExt_uid88_fpAddTest_q_a8_a.is_wysiwyg = "true";
defparam fp_functions_0_aleftShiftStage2_uid249_fracPostNormExt_uid88_fpAddTest_q_a8_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aleftShiftStage2_uid249_fracPostNormExt_uid88_fpAddTest_q_a9_a(
	.clk(clk),
	.d(fp_functions_0_ai3365_a4_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aleftShiftStage2_uid249_fracPostNormExt_uid88_fpAddTest_q_a9_a_aq));
defparam fp_functions_0_aleftShiftStage2_uid249_fracPostNormExt_uid88_fpAddTest_q_a9_a.is_wysiwyg = "true";
defparam fp_functions_0_aleftShiftStage2_uid249_fracPostNormExt_uid88_fpAddTest_q_a9_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aleftShiftStage2_uid249_fracPostNormExt_uid88_fpAddTest_q_a10_a(
	.clk(clk),
	.d(fp_functions_0_ai3365_a5_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aleftShiftStage2_uid249_fracPostNormExt_uid88_fpAddTest_q_a10_a_aq));
defparam fp_functions_0_aleftShiftStage2_uid249_fracPostNormExt_uid88_fpAddTest_q_a10_a.is_wysiwyg = "true";
defparam fp_functions_0_aleftShiftStage2_uid249_fracPostNormExt_uid88_fpAddTest_q_a10_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aleftShiftStage2_uid249_fracPostNormExt_uid88_fpAddTest_q_a11_a(
	.clk(clk),
	.d(fp_functions_0_ai3365_a6_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aleftShiftStage2_uid249_fracPostNormExt_uid88_fpAddTest_q_a11_a_aq));
defparam fp_functions_0_aleftShiftStage2_uid249_fracPostNormExt_uid88_fpAddTest_q_a11_a.is_wysiwyg = "true";
defparam fp_functions_0_aleftShiftStage2_uid249_fracPostNormExt_uid88_fpAddTest_q_a11_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aleftShiftStage2_uid249_fracPostNormExt_uid88_fpAddTest_q_a12_a(
	.clk(clk),
	.d(fp_functions_0_ai3365_a7_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aleftShiftStage2_uid249_fracPostNormExt_uid88_fpAddTest_q_a12_a_aq));
defparam fp_functions_0_aleftShiftStage2_uid249_fracPostNormExt_uid88_fpAddTest_q_a12_a.is_wysiwyg = "true";
defparam fp_functions_0_aleftShiftStage2_uid249_fracPostNormExt_uid88_fpAddTest_q_a12_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aleftShiftStage2_uid249_fracPostNormExt_uid88_fpAddTest_q_a13_a(
	.clk(clk),
	.d(fp_functions_0_ai3365_a8_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aleftShiftStage2_uid249_fracPostNormExt_uid88_fpAddTest_q_a13_a_aq));
defparam fp_functions_0_aleftShiftStage2_uid249_fracPostNormExt_uid88_fpAddTest_q_a13_a.is_wysiwyg = "true";
defparam fp_functions_0_aleftShiftStage2_uid249_fracPostNormExt_uid88_fpAddTest_q_a13_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aleftShiftStage2_uid249_fracPostNormExt_uid88_fpAddTest_q_a14_a(
	.clk(clk),
	.d(fp_functions_0_ai3365_a9_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aleftShiftStage2_uid249_fracPostNormExt_uid88_fpAddTest_q_a14_a_aq));
defparam fp_functions_0_aleftShiftStage2_uid249_fracPostNormExt_uid88_fpAddTest_q_a14_a.is_wysiwyg = "true";
defparam fp_functions_0_aleftShiftStage2_uid249_fracPostNormExt_uid88_fpAddTest_q_a14_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aleftShiftStage2_uid249_fracPostNormExt_uid88_fpAddTest_q_a15_a(
	.clk(clk),
	.d(fp_functions_0_ai3365_a10_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aleftShiftStage2_uid249_fracPostNormExt_uid88_fpAddTest_q_a15_a_aq));
defparam fp_functions_0_aleftShiftStage2_uid249_fracPostNormExt_uid88_fpAddTest_q_a15_a.is_wysiwyg = "true";
defparam fp_functions_0_aleftShiftStage2_uid249_fracPostNormExt_uid88_fpAddTest_q_a15_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aleftShiftStage2_uid249_fracPostNormExt_uid88_fpAddTest_q_a16_a(
	.clk(clk),
	.d(fp_functions_0_ai3365_a11_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aleftShiftStage2_uid249_fracPostNormExt_uid88_fpAddTest_q_a16_a_aq));
defparam fp_functions_0_aleftShiftStage2_uid249_fracPostNormExt_uid88_fpAddTest_q_a16_a.is_wysiwyg = "true";
defparam fp_functions_0_aleftShiftStage2_uid249_fracPostNormExt_uid88_fpAddTest_q_a16_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aleftShiftStage2_uid249_fracPostNormExt_uid88_fpAddTest_q_a17_a(
	.clk(clk),
	.d(fp_functions_0_ai3365_a12_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aleftShiftStage2_uid249_fracPostNormExt_uid88_fpAddTest_q_a17_a_aq));
defparam fp_functions_0_aleftShiftStage2_uid249_fracPostNormExt_uid88_fpAddTest_q_a17_a.is_wysiwyg = "true";
defparam fp_functions_0_aleftShiftStage2_uid249_fracPostNormExt_uid88_fpAddTest_q_a17_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aleftShiftStage2_uid249_fracPostNormExt_uid88_fpAddTest_q_a18_a(
	.clk(clk),
	.d(fp_functions_0_ai3365_a13_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aleftShiftStage2_uid249_fracPostNormExt_uid88_fpAddTest_q_a18_a_aq));
defparam fp_functions_0_aleftShiftStage2_uid249_fracPostNormExt_uid88_fpAddTest_q_a18_a.is_wysiwyg = "true";
defparam fp_functions_0_aleftShiftStage2_uid249_fracPostNormExt_uid88_fpAddTest_q_a18_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aleftShiftStage2_uid249_fracPostNormExt_uid88_fpAddTest_q_a19_a(
	.clk(clk),
	.d(fp_functions_0_ai3365_a14_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aleftShiftStage2_uid249_fracPostNormExt_uid88_fpAddTest_q_a19_a_aq));
defparam fp_functions_0_aleftShiftStage2_uid249_fracPostNormExt_uid88_fpAddTest_q_a19_a.is_wysiwyg = "true";
defparam fp_functions_0_aleftShiftStage2_uid249_fracPostNormExt_uid88_fpAddTest_q_a19_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aleftShiftStage2_uid249_fracPostNormExt_uid88_fpAddTest_q_a20_a(
	.clk(clk),
	.d(fp_functions_0_ai3365_a15_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aleftShiftStage2_uid249_fracPostNormExt_uid88_fpAddTest_q_a20_a_aq));
defparam fp_functions_0_aleftShiftStage2_uid249_fracPostNormExt_uid88_fpAddTest_q_a20_a.is_wysiwyg = "true";
defparam fp_functions_0_aleftShiftStage2_uid249_fracPostNormExt_uid88_fpAddTest_q_a20_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aleftShiftStage2_uid249_fracPostNormExt_uid88_fpAddTest_q_a21_a(
	.clk(clk),
	.d(fp_functions_0_ai3365_a16_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aleftShiftStage2_uid249_fracPostNormExt_uid88_fpAddTest_q_a21_a_aq));
defparam fp_functions_0_aleftShiftStage2_uid249_fracPostNormExt_uid88_fpAddTest_q_a21_a.is_wysiwyg = "true";
defparam fp_functions_0_aleftShiftStage2_uid249_fracPostNormExt_uid88_fpAddTest_q_a21_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aleftShiftStage2_uid249_fracPostNormExt_uid88_fpAddTest_q_a22_a(
	.clk(clk),
	.d(fp_functions_0_ai3365_a17_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aleftShiftStage2_uid249_fracPostNormExt_uid88_fpAddTest_q_a22_a_aq));
defparam fp_functions_0_aleftShiftStage2_uid249_fracPostNormExt_uid88_fpAddTest_q_a22_a.is_wysiwyg = "true";
defparam fp_functions_0_aleftShiftStage2_uid249_fracPostNormExt_uid88_fpAddTest_q_a22_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aleftShiftStage2_uid249_fracPostNormExt_uid88_fpAddTest_q_a23_a(
	.clk(clk),
	.d(fp_functions_0_ai3337_a1_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aleftShiftStage2_uid249_fracPostNormExt_uid88_fpAddTest_q_a23_a_aq));
defparam fp_functions_0_aleftShiftStage2_uid249_fracPostNormExt_uid88_fpAddTest_q_a23_a.is_wysiwyg = "true";
defparam fp_functions_0_aleftShiftStage2_uid249_fracPostNormExt_uid88_fpAddTest_q_a23_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aleftShiftStage2_uid249_fracPostNormExt_uid88_fpAddTest_q_a24_a(
	.clk(clk),
	.d(fp_functions_0_ai3365_a18_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aleftShiftStage2_uid249_fracPostNormExt_uid88_fpAddTest_q_a24_a_aq));
defparam fp_functions_0_aleftShiftStage2_uid249_fracPostNormExt_uid88_fpAddTest_q_a24_a.is_wysiwyg = "true";
defparam fp_functions_0_aleftShiftStage2_uid249_fracPostNormExt_uid88_fpAddTest_q_a24_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aleftShiftStage2_uid249_fracPostNormExt_uid88_fpAddTest_q_a25_a(
	.clk(clk),
	.d(fp_functions_0_ai3365_a19_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aleftShiftStage2_uid249_fracPostNormExt_uid88_fpAddTest_q_a25_a_aq));
defparam fp_functions_0_aleftShiftStage2_uid249_fracPostNormExt_uid88_fpAddTest_q_a25_a.is_wysiwyg = "true";
defparam fp_functions_0_aleftShiftStage2_uid249_fracPostNormExt_uid88_fpAddTest_q_a25_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aleftShiftStage2_uid249_fracPostNormExt_uid88_fpAddTest_q_a26_a(
	.clk(clk),
	.d(fp_functions_0_ai3337_a2_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aleftShiftStage2_uid249_fracPostNormExt_uid88_fpAddTest_q_a26_a_aq));
defparam fp_functions_0_aleftShiftStage2_uid249_fracPostNormExt_uid88_fpAddTest_q_a26_a.is_wysiwyg = "true";
defparam fp_functions_0_aleftShiftStage2_uid249_fracPostNormExt_uid88_fpAddTest_q_a26_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist6_sigB_uid51_fpAddTest_b_2_q_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist5_sigB_uid51_fpAddTest_b_1_q_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist6_sigB_uid51_fpAddTest_b_2_q_a0_a_aq));
defparam fp_functions_0_aredist6_sigB_uid51_fpAddTest_b_2_q_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist6_sigB_uid51_fpAddTest_b_2_q_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist8_sigA_uid50_fpAddTest_b_2_q_a0_a(
	.clk(clk),
	.d(fp_functions_0_aredist7_sigA_uid50_fpAddTest_b_1_q_a0_a_aq),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist8_sigA_uid50_fpAddTest_b_2_q_a0_a_aq));
defparam fp_functions_0_aredist8_sigA_uid50_fpAddTest_b_2_q_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist8_sigA_uid50_fpAddTest_b_2_q_a0_a.power_up = "dont_care";

fourteennm_lcell_comb fp_functions_0_aadd_4_a1(
	.dataa(!fp_functions_0_aredist7_sigA_uid50_fpAddTest_b_1_q_a0_a_aq),
	.datab(!fp_functions_0_aredist5_sigB_uid51_fpAddTest_b_1_q_a0_a_aq),
	.datac(!fp_functions_0_aredist17_frac_aSig_uid22_fpAddTest_b_1_q_a17_a_aq),
	.datad(!fp_functions_0_astickyBits_uid69_fpAddTest_merged_bit_select_b_a0_a_a0_combout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_4_a42),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_4_a1_sumout),
	.cout(fp_functions_0_aadd_4_a2),
	.shareout());
defparam fp_functions_0_aadd_4_a1.extended_lut = "off";
defparam fp_functions_0_aadd_4_a1.lut_mask = 64'h0000000006096996;
defparam fp_functions_0_aadd_4_a1.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_4_a6(
	.dataa(!fp_functions_0_aredist7_sigA_uid50_fpAddTest_b_1_q_a0_a_aq),
	.datab(!fp_functions_0_aredist5_sigB_uid51_fpAddTest_b_1_q_a0_a_aq),
	.datac(!fp_functions_0_aredist17_frac_aSig_uid22_fpAddTest_b_1_q_a13_a_aq),
	.datad(!fp_functions_0_astickyBits_uid69_fpAddTest_merged_bit_select_b_a0_a_a1_combout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_4_a27),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_4_a6_sumout),
	.cout(fp_functions_0_aadd_4_a7),
	.shareout());
defparam fp_functions_0_aadd_4_a6.extended_lut = "off";
defparam fp_functions_0_aadd_4_a6.lut_mask = 64'h0000000006096996;
defparam fp_functions_0_aadd_4_a6.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_4_a11(
	.dataa(!fp_functions_0_aredist7_sigA_uid50_fpAddTest_b_1_q_a0_a_aq),
	.datab(!fp_functions_0_aredist5_sigB_uid51_fpAddTest_b_1_q_a0_a_aq),
	.datac(!fp_functions_0_aredist17_frac_aSig_uid22_fpAddTest_b_1_q_a9_a_aq),
	.datad(!fp_functions_0_astickyBits_uid69_fpAddTest_merged_bit_select_b_a0_a_a2_combout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_4_a102),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_4_a11_sumout),
	.cout(fp_functions_0_aadd_4_a12),
	.shareout());
defparam fp_functions_0_aadd_4_a11.extended_lut = "off";
defparam fp_functions_0_aadd_4_a11.lut_mask = 64'h0000000006096996;
defparam fp_functions_0_aadd_4_a11.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_4_a16(
	.dataa(!fp_functions_0_aredist7_sigA_uid50_fpAddTest_b_1_q_a0_a_aq),
	.datab(!fp_functions_0_aredist5_sigB_uid51_fpAddTest_b_1_q_a0_a_aq),
	.datac(!fp_functions_0_aredist17_frac_aSig_uid22_fpAddTest_b_1_q_a10_a_aq),
	.datad(!fp_functions_0_astickyBits_uid69_fpAddTest_merged_bit_select_b_a0_a_a3_combout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_4_a12),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_4_a16_sumout),
	.cout(fp_functions_0_aadd_4_a17),
	.shareout());
defparam fp_functions_0_aadd_4_a16.extended_lut = "off";
defparam fp_functions_0_aadd_4_a16.lut_mask = 64'h0000000006096996;
defparam fp_functions_0_aadd_4_a16.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_4_a21(
	.dataa(!fp_functions_0_aredist7_sigA_uid50_fpAddTest_b_1_q_a0_a_aq),
	.datab(!fp_functions_0_aredist5_sigB_uid51_fpAddTest_b_1_q_a0_a_aq),
	.datac(!fp_functions_0_aredist17_frac_aSig_uid22_fpAddTest_b_1_q_a11_a_aq),
	.datad(!fp_functions_0_astickyBits_uid69_fpAddTest_merged_bit_select_b_a0_a_a4_combout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_4_a17),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_4_a21_sumout),
	.cout(fp_functions_0_aadd_4_a22),
	.shareout());
defparam fp_functions_0_aadd_4_a21.extended_lut = "off";
defparam fp_functions_0_aadd_4_a21.lut_mask = 64'h0000000006096996;
defparam fp_functions_0_aadd_4_a21.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_4_a26(
	.dataa(!fp_functions_0_aredist7_sigA_uid50_fpAddTest_b_1_q_a0_a_aq),
	.datab(!fp_functions_0_aredist5_sigB_uid51_fpAddTest_b_1_q_a0_a_aq),
	.datac(!fp_functions_0_aredist17_frac_aSig_uid22_fpAddTest_b_1_q_a12_a_aq),
	.datad(!fp_functions_0_astickyBits_uid69_fpAddTest_merged_bit_select_b_a0_a_a5_combout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_4_a22),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_4_a26_sumout),
	.cout(fp_functions_0_aadd_4_a27),
	.shareout());
defparam fp_functions_0_aadd_4_a26.extended_lut = "off";
defparam fp_functions_0_aadd_4_a26.lut_mask = 64'h0000000006096996;
defparam fp_functions_0_aadd_4_a26.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_4_a31(
	.dataa(!fp_functions_0_aredist7_sigA_uid50_fpAddTest_b_1_q_a0_a_aq),
	.datab(!fp_functions_0_aredist5_sigB_uid51_fpAddTest_b_1_q_a0_a_aq),
	.datac(!fp_functions_0_aredist17_frac_aSig_uid22_fpAddTest_b_1_q_a14_a_aq),
	.datad(!fp_functions_0_astickyBits_uid69_fpAddTest_merged_bit_select_b_a0_a_a6_combout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_4_a7),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_4_a31_sumout),
	.cout(fp_functions_0_aadd_4_a32),
	.shareout());
defparam fp_functions_0_aadd_4_a31.extended_lut = "off";
defparam fp_functions_0_aadd_4_a31.lut_mask = 64'h0000000006096996;
defparam fp_functions_0_aadd_4_a31.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_4_a36(
	.dataa(!fp_functions_0_aredist7_sigA_uid50_fpAddTest_b_1_q_a0_a_aq),
	.datab(!fp_functions_0_aredist5_sigB_uid51_fpAddTest_b_1_q_a0_a_aq),
	.datac(!fp_functions_0_aredist17_frac_aSig_uid22_fpAddTest_b_1_q_a15_a_aq),
	.datad(!fp_functions_0_astickyBits_uid69_fpAddTest_merged_bit_select_b_a0_a_a7_combout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_4_a32),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_4_a36_sumout),
	.cout(fp_functions_0_aadd_4_a37),
	.shareout());
defparam fp_functions_0_aadd_4_a36.extended_lut = "off";
defparam fp_functions_0_aadd_4_a36.lut_mask = 64'h0000000006096996;
defparam fp_functions_0_aadd_4_a36.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_4_a41(
	.dataa(!fp_functions_0_aredist7_sigA_uid50_fpAddTest_b_1_q_a0_a_aq),
	.datab(!fp_functions_0_aredist5_sigB_uid51_fpAddTest_b_1_q_a0_a_aq),
	.datac(!fp_functions_0_aredist17_frac_aSig_uid22_fpAddTest_b_1_q_a16_a_aq),
	.datad(!fp_functions_0_astickyBits_uid69_fpAddTest_merged_bit_select_b_a0_a_a8_combout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_4_a37),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_4_a41_sumout),
	.cout(fp_functions_0_aadd_4_a42),
	.shareout());
defparam fp_functions_0_aadd_4_a41.extended_lut = "off";
defparam fp_functions_0_aadd_4_a41.lut_mask = 64'h0000000006096996;
defparam fp_functions_0_aadd_4_a41.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_4_a46(
	.dataa(!fp_functions_0_aredist5_sigB_uid51_fpAddTest_b_1_q_a0_a_aq),
	.datab(!fp_functions_0_aredist7_sigA_uid50_fpAddTest_b_1_q_a0_a_aq),
	.datac(!fp_functions_0_aredist17_frac_aSig_uid22_fpAddTest_b_1_q_a22_a_aq),
	.datad(!fp_functions_0_astickyBits_uid69_fpAddTest_merged_bit_select_b_a0_a_a9_combout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_4_a72),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_4_a46_sumout),
	.cout(fp_functions_0_aadd_4_a47),
	.shareout());
defparam fp_functions_0_aadd_4_a46.extended_lut = "off";
defparam fp_functions_0_aadd_4_a46.lut_mask = 64'h0000000006096996;
defparam fp_functions_0_aadd_4_a46.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_4_a51(
	.dataa(!fp_functions_0_aredist5_sigB_uid51_fpAddTest_b_1_q_a0_a_aq),
	.datab(!fp_functions_0_aredist7_sigA_uid50_fpAddTest_b_1_q_a0_a_aq),
	.datac(!fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a48_a_aq),
	.datad(!fp_functions_0_ashiftedOut_uid63_fpAddTest_o_a10_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_4_a47),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_4_a51_sumout),
	.cout(fp_functions_0_aadd_4_a52),
	.shareout());
defparam fp_functions_0_aadd_4_a51.extended_lut = "off";
defparam fp_functions_0_aadd_4_a51.lut_mask = 64'h0000000069669699;
defparam fp_functions_0_aadd_4_a51.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_4_a56(
	.dataa(!fp_functions_0_aredist7_sigA_uid50_fpAddTest_b_1_q_a0_a_aq),
	.datab(!fp_functions_0_aredist5_sigB_uid51_fpAddTest_b_1_q_a0_a_aq),
	.datac(!fp_functions_0_aredist17_frac_aSig_uid22_fpAddTest_b_1_q_a18_a_aq),
	.datad(!fp_functions_0_astickyBits_uid69_fpAddTest_merged_bit_select_b_a0_a_a10_combout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_4_a2),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_4_a56_sumout),
	.cout(fp_functions_0_aadd_4_a57),
	.shareout());
defparam fp_functions_0_aadd_4_a56.extended_lut = "off";
defparam fp_functions_0_aadd_4_a56.lut_mask = 64'h0000000006096996;
defparam fp_functions_0_aadd_4_a56.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_4_a61(
	.dataa(!fp_functions_0_aredist7_sigA_uid50_fpAddTest_b_1_q_a0_a_aq),
	.datab(!fp_functions_0_aredist5_sigB_uid51_fpAddTest_b_1_q_a0_a_aq),
	.datac(!fp_functions_0_aredist17_frac_aSig_uid22_fpAddTest_b_1_q_a19_a_aq),
	.datad(!fp_functions_0_astickyBits_uid69_fpAddTest_merged_bit_select_b_a0_a_a11_combout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_4_a57),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_4_a61_sumout),
	.cout(fp_functions_0_aadd_4_a62),
	.shareout());
defparam fp_functions_0_aadd_4_a61.extended_lut = "off";
defparam fp_functions_0_aadd_4_a61.lut_mask = 64'h0000000006096996;
defparam fp_functions_0_aadd_4_a61.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_4_a66(
	.dataa(!fp_functions_0_aredist7_sigA_uid50_fpAddTest_b_1_q_a0_a_aq),
	.datab(!fp_functions_0_aredist5_sigB_uid51_fpAddTest_b_1_q_a0_a_aq),
	.datac(!fp_functions_0_aredist17_frac_aSig_uid22_fpAddTest_b_1_q_a20_a_aq),
	.datad(!fp_functions_0_astickyBits_uid69_fpAddTest_merged_bit_select_b_a0_a_a12_combout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_4_a62),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_4_a66_sumout),
	.cout(fp_functions_0_aadd_4_a67),
	.shareout());
defparam fp_functions_0_aadd_4_a66.extended_lut = "off";
defparam fp_functions_0_aadd_4_a66.lut_mask = 64'h0000000006096996;
defparam fp_functions_0_aadd_4_a66.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_4_a71(
	.dataa(!fp_functions_0_aredist7_sigA_uid50_fpAddTest_b_1_q_a0_a_aq),
	.datab(!fp_functions_0_aredist5_sigB_uid51_fpAddTest_b_1_q_a0_a_aq),
	.datac(!fp_functions_0_aredist17_frac_aSig_uid22_fpAddTest_b_1_q_a21_a_aq),
	.datad(!fp_functions_0_astickyBits_uid69_fpAddTest_merged_bit_select_b_a0_a_a13_combout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_4_a67),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_4_a71_sumout),
	.cout(fp_functions_0_aadd_4_a72),
	.shareout());
defparam fp_functions_0_aadd_4_a71.extended_lut = "off";
defparam fp_functions_0_aadd_4_a71.lut_mask = 64'h0000000006096996;
defparam fp_functions_0_aadd_4_a71.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_4_a76(
	.dataa(!fp_functions_0_aredist5_sigB_uid51_fpAddTest_b_1_q_a0_a_aq),
	.datab(gnd),
	.datac(!fp_functions_0_aredist7_sigA_uid50_fpAddTest_b_1_q_a0_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_4_a52),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_4_a76_sumout),
	.cout(),
	.shareout());
defparam fp_functions_0_aadd_4_a76.extended_lut = "off";
defparam fp_functions_0_aadd_4_a76.lut_mask = 64'h0000000000005A5A;
defparam fp_functions_0_aadd_4_a76.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_4_a81(
	.dataa(!fp_functions_0_aredist7_sigA_uid50_fpAddTest_b_1_q_a0_a_aq),
	.datab(!fp_functions_0_aredist5_sigB_uid51_fpAddTest_b_1_q_a0_a_aq),
	.datac(!fp_functions_0_aredist17_frac_aSig_uid22_fpAddTest_b_1_q_a4_a_aq),
	.datad(!fp_functions_0_astickyBits_uid69_fpAddTest_merged_bit_select_b_a0_a_a14_combout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_4_a87),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_4_a81_sumout),
	.cout(fp_functions_0_aadd_4_a82),
	.shareout());
defparam fp_functions_0_aadd_4_a81.extended_lut = "off";
defparam fp_functions_0_aadd_4_a81.lut_mask = 64'h0000000006096996;
defparam fp_functions_0_aadd_4_a81.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_4_a86(
	.dataa(!fp_functions_0_aredist7_sigA_uid50_fpAddTest_b_1_q_a0_a_aq),
	.datab(!fp_functions_0_aredist5_sigB_uid51_fpAddTest_b_1_q_a0_a_aq),
	.datac(!fp_functions_0_aredist17_frac_aSig_uid22_fpAddTest_b_1_q_a3_a_aq),
	.datad(!fp_functions_0_astickyBits_uid69_fpAddTest_merged_bit_select_b_a0_a_a15_combout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_4_a97),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_4_a86_sumout),
	.cout(fp_functions_0_aadd_4_a87),
	.shareout());
defparam fp_functions_0_aadd_4_a86.extended_lut = "off";
defparam fp_functions_0_aadd_4_a86.lut_mask = 64'h0000000006096996;
defparam fp_functions_0_aadd_4_a86.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_4_a91(
	.dataa(!fp_functions_0_aredist7_sigA_uid50_fpAddTest_b_1_q_a0_a_aq),
	.datab(!fp_functions_0_aredist5_sigB_uid51_fpAddTest_b_1_q_a0_a_aq),
	.datac(!fp_functions_0_aredist17_frac_aSig_uid22_fpAddTest_b_1_q_a1_a_aq),
	.datad(!fp_functions_0_astickyBits_uid69_fpAddTest_merged_bit_select_b_a0_a_a16_combout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_4_a112),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_4_a91_sumout),
	.cout(fp_functions_0_aadd_4_a92),
	.shareout());
defparam fp_functions_0_aadd_4_a91.extended_lut = "off";
defparam fp_functions_0_aadd_4_a91.lut_mask = 64'h0000000006096996;
defparam fp_functions_0_aadd_4_a91.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_4_a96(
	.dataa(!fp_functions_0_aredist7_sigA_uid50_fpAddTest_b_1_q_a0_a_aq),
	.datab(!fp_functions_0_aredist5_sigB_uid51_fpAddTest_b_1_q_a0_a_aq),
	.datac(!fp_functions_0_aredist17_frac_aSig_uid22_fpAddTest_b_1_q_a2_a_aq),
	.datad(!fp_functions_0_astickyBits_uid69_fpAddTest_merged_bit_select_b_a0_a_a17_combout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_4_a92),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_4_a96_sumout),
	.cout(fp_functions_0_aadd_4_a97),
	.shareout());
defparam fp_functions_0_aadd_4_a96.extended_lut = "off";
defparam fp_functions_0_aadd_4_a96.lut_mask = 64'h0000000006096996;
defparam fp_functions_0_aadd_4_a96.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_4_a101(
	.dataa(!fp_functions_0_aredist7_sigA_uid50_fpAddTest_b_1_q_a0_a_aq),
	.datab(!fp_functions_0_aredist5_sigB_uid51_fpAddTest_b_1_q_a0_a_aq),
	.datac(!fp_functions_0_aredist17_frac_aSig_uid22_fpAddTest_b_1_q_a8_a_aq),
	.datad(!fp_functions_0_astickyBits_uid69_fpAddTest_merged_bit_select_b_a0_a_a18_combout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_4_a107),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_4_a101_sumout),
	.cout(fp_functions_0_aadd_4_a102),
	.shareout());
defparam fp_functions_0_aadd_4_a101.extended_lut = "off";
defparam fp_functions_0_aadd_4_a101.lut_mask = 64'h0000000006096996;
defparam fp_functions_0_aadd_4_a101.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_4_a106(
	.dataa(!fp_functions_0_aredist7_sigA_uid50_fpAddTest_b_1_q_a0_a_aq),
	.datab(!fp_functions_0_aredist5_sigB_uid51_fpAddTest_b_1_q_a0_a_aq),
	.datac(!fp_functions_0_aredist17_frac_aSig_uid22_fpAddTest_b_1_q_a7_a_aq),
	.datad(!fp_functions_0_astickyBits_uid69_fpAddTest_merged_bit_select_b_a0_a_a19_combout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_4_a122),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_4_a106_sumout),
	.cout(fp_functions_0_aadd_4_a107),
	.shareout());
defparam fp_functions_0_aadd_4_a106.extended_lut = "off";
defparam fp_functions_0_aadd_4_a106.lut_mask = 64'h0000000006096996;
defparam fp_functions_0_aadd_4_a106.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_4_a111(
	.dataa(!fp_functions_0_aredist7_sigA_uid50_fpAddTest_b_1_q_a0_a_aq),
	.datab(!fp_functions_0_aredist5_sigB_uid51_fpAddTest_b_1_q_a0_a_aq),
	.datac(!fp_functions_0_aredist17_frac_aSig_uid22_fpAddTest_b_1_q_a0_a_aq),
	.datad(!fp_functions_0_astickyBits_uid69_fpAddTest_merged_bit_select_b_a0_a_a20_combout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_4_a127),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_4_a111_sumout),
	.cout(fp_functions_0_aadd_4_a112),
	.shareout());
defparam fp_functions_0_aadd_4_a111.extended_lut = "off";
defparam fp_functions_0_aadd_4_a111.lut_mask = 64'h0000000006096996;
defparam fp_functions_0_aadd_4_a111.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_4_a116(
	.dataa(!fp_functions_0_aredist7_sigA_uid50_fpAddTest_b_1_q_a0_a_aq),
	.datab(!fp_functions_0_aredist5_sigB_uid51_fpAddTest_b_1_q_a0_a_aq),
	.datac(!fp_functions_0_aredist17_frac_aSig_uid22_fpAddTest_b_1_q_a5_a_aq),
	.datad(!fp_functions_0_astickyBits_uid69_fpAddTest_merged_bit_select_b_a0_a_a21_combout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_4_a82),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_4_a116_sumout),
	.cout(fp_functions_0_aadd_4_a117),
	.shareout());
defparam fp_functions_0_aadd_4_a116.extended_lut = "off";
defparam fp_functions_0_aadd_4_a116.lut_mask = 64'h0000000006096996;
defparam fp_functions_0_aadd_4_a116.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_4_a121(
	.dataa(!fp_functions_0_aredist7_sigA_uid50_fpAddTest_b_1_q_a0_a_aq),
	.datab(!fp_functions_0_aredist5_sigB_uid51_fpAddTest_b_1_q_a0_a_aq),
	.datac(!fp_functions_0_aredist17_frac_aSig_uid22_fpAddTest_b_1_q_a6_a_aq),
	.datad(!fp_functions_0_astickyBits_uid69_fpAddTest_merged_bit_select_b_a0_a_a22_combout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_4_a117),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_4_a121_sumout),
	.cout(fp_functions_0_aadd_4_a122),
	.shareout());
defparam fp_functions_0_aadd_4_a121.extended_lut = "off";
defparam fp_functions_0_aadd_4_a121.lut_mask = 64'h0000000006096996;
defparam fp_functions_0_aadd_4_a121.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_4_a126(
	.dataa(!fp_functions_0_aredist5_sigB_uid51_fpAddTest_b_1_q_a0_a_aq),
	.datab(!fp_functions_0_aredist7_sigA_uid50_fpAddTest_b_1_q_a0_a_aq),
	.datac(!fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a24_a_aq),
	.datad(!fp_functions_0_ashiftedOut_uid63_fpAddTest_o_a10_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_4_a132),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_4_a126_sumout),
	.cout(fp_functions_0_aadd_4_a127),
	.shareout());
defparam fp_functions_0_aadd_4_a126.extended_lut = "off";
defparam fp_functions_0_aadd_4_a126.lut_mask = 64'h0000000000006966;
defparam fp_functions_0_aadd_4_a126.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_4_a131(
	.dataa(!fp_functions_0_aredist5_sigB_uid51_fpAddTest_b_1_q_a0_a_aq),
	.datab(!fp_functions_0_aredist7_sigA_uid50_fpAddTest_b_1_q_a0_a_aq),
	.datac(!fp_functions_0_areduce_nor_1_a4_combout),
	.datad(!fp_functions_0_astickyBits_uid69_fpAddTest_merged_bit_select_b_a0_a_a23_combout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_4_a131_sumout),
	.cout(fp_functions_0_aadd_4_a132),
	.shareout());
defparam fp_functions_0_aadd_4_a131.extended_lut = "off";
defparam fp_functions_0_aadd_4_a131.lut_mask = 64'h00000000600006F9;
defparam fp_functions_0_aadd_4_a131.shared_arith = "off";

fourteennm_ff fp_functions_0_ashiftedOut_uid63_fpAddTest_o_a10_a(
	.clk(clk),
	.d(fp_functions_0_aadd_2_a1_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_ashiftedOut_uid63_fpAddTest_o_a10_a_aq));
defparam fp_functions_0_ashiftedOut_uid63_fpAddTest_o_a10_a.is_wysiwyg = "true";
defparam fp_functions_0_ashiftedOut_uid63_fpAddTest_o_a10_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a22_a(
	.clk(clk),
	.d(fp_functions_0_ai1783_a0_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a28_a_a0_combout),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a22_a_aq));
defparam fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a22_a.is_wysiwyg = "true";
defparam fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a22_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a16_a(
	.clk(clk),
	.d(fp_functions_0_ai1734_a1_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a16_a_aq));
defparam fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a16_a.is_wysiwyg = "true";
defparam fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a16_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a0_a(
	.clk(clk),
	.d(fp_functions_0_ai1734_a2_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a0_a_aq));
defparam fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a1_a(
	.clk(clk),
	.d(fp_functions_0_ai1783_a1_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a2_a_a1_combout),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a1_a_aq));
defparam fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a1_a.is_wysiwyg = "true";
defparam fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a1_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a9_a(
	.clk(clk),
	.d(fp_functions_0_ai1783_a2_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a2_a_a1_combout),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a9_a_aq));
defparam fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a9_a.is_wysiwyg = "true";
defparam fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a9_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a4_a(
	.clk(clk),
	.d(fp_functions_0_ai1783_a3_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a2_a_a1_combout),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a4_a_aq));
defparam fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a4_a.is_wysiwyg = "true";
defparam fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a4_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a21_a(
	.clk(clk),
	.d(fp_functions_0_ai1783_a4_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a28_a_a0_combout),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a21_a_aq));
defparam fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a21_a.is_wysiwyg = "true";
defparam fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a21_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a20_a(
	.clk(clk),
	.d(fp_functions_0_ai1783_a5_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a28_a_a0_combout),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a20_a_aq));
defparam fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a20_a.is_wysiwyg = "true";
defparam fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a20_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a19_a(
	.clk(clk),
	.d(fp_functions_0_ai1783_a6_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a28_a_a0_combout),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a19_a_aq));
defparam fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a19_a.is_wysiwyg = "true";
defparam fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a19_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a17_a(
	.clk(clk),
	.d(fp_functions_0_ai1783_a7_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a28_a_a0_combout),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a17_a_aq));
defparam fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a17_a.is_wysiwyg = "true";
defparam fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a17_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a18_a(
	.clk(clk),
	.d(fp_functions_0_ai1783_a8_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a28_a_a0_combout),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a18_a_aq));
defparam fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a18_a.is_wysiwyg = "true";
defparam fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a18_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a8_a(
	.clk(clk),
	.d(fp_functions_0_ai1783_a9_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a2_a_a1_combout),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a8_a_aq));
defparam fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a8_a.is_wysiwyg = "true";
defparam fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a8_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a7_a(
	.clk(clk),
	.d(fp_functions_0_ai1783_a11_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a2_a_a1_combout),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a7_a_aq));
defparam fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a7_a.is_wysiwyg = "true";
defparam fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a7_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a6_a(
	.clk(clk),
	.d(fp_functions_0_ai1783_a12_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a2_a_a1_combout),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a6_a_aq));
defparam fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a6_a.is_wysiwyg = "true";
defparam fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a6_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a5_a(
	.clk(clk),
	.d(fp_functions_0_ai1783_a13_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a2_a_a1_combout),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a5_a_aq));
defparam fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a5_a.is_wysiwyg = "true";
defparam fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a5_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a2_a(
	.clk(clk),
	.d(fp_functions_0_ai1783_a14_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a2_a_a1_combout),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a2_a_aq));
defparam fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a2_a.is_wysiwyg = "true";
defparam fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a2_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a3_a(
	.clk(clk),
	.d(fp_functions_0_ai1783_a15_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a2_a_a1_combout),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a3_a_aq));
defparam fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a3_a.is_wysiwyg = "true";
defparam fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a3_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aexpXIsMax_uid38_fpAddTest_delay_adelay_signals_a0_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_areduce_nor_7_a3_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aexpXIsMax_uid38_fpAddTest_delay_adelay_signals_a0_a_a0_a_aq));
defparam fp_functions_0_aexpXIsMax_uid38_fpAddTest_delay_adelay_signals_a0_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aexpXIsMax_uid38_fpAddTest_delay_adelay_signals_a0_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist9_InvExpXIsZero_uid44_fpAddTest_q_2_delay_0_a0_a(
	.clk(clk),
	.d(fp_functions_0_areduce_nor_0_acombout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist9_InvExpXIsZero_uid44_fpAddTest_q_2_delay_0_a0_a_aq));
defparam fp_functions_0_aredist9_InvExpXIsZero_uid44_fpAddTest_q_2_delay_0_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist9_InvExpXIsZero_uid44_fpAddTest_q_2_delay_0_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist18_exp_aSig_uid21_fpAddTest_b_2_delay_0_a4_a(
	.clk(clk),
	.d(fp_functions_0_aexp_aSig_uid21_fpAddTest_b_a0_a_a0_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist18_exp_aSig_uid21_fpAddTest_b_2_delay_0_a4_a_aq));
defparam fp_functions_0_aredist18_exp_aSig_uid21_fpAddTest_b_2_delay_0_a4_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist18_exp_aSig_uid21_fpAddTest_b_2_delay_0_a4_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist18_exp_aSig_uid21_fpAddTest_b_2_delay_0_a5_a(
	.clk(clk),
	.d(fp_functions_0_aexp_aSig_uid21_fpAddTest_b_a0_a_a1_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist18_exp_aSig_uid21_fpAddTest_b_2_delay_0_a5_a_aq));
defparam fp_functions_0_aredist18_exp_aSig_uid21_fpAddTest_b_2_delay_0_a5_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist18_exp_aSig_uid21_fpAddTest_b_2_delay_0_a5_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist18_exp_aSig_uid21_fpAddTest_b_2_delay_0_a6_a(
	.clk(clk),
	.d(fp_functions_0_aexp_aSig_uid21_fpAddTest_b_a0_a_a2_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist18_exp_aSig_uid21_fpAddTest_b_2_delay_0_a6_a_aq));
defparam fp_functions_0_aredist18_exp_aSig_uid21_fpAddTest_b_2_delay_0_a6_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist18_exp_aSig_uid21_fpAddTest_b_2_delay_0_a6_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist18_exp_aSig_uid21_fpAddTest_b_2_delay_0_a7_a(
	.clk(clk),
	.d(fp_functions_0_aexp_aSig_uid21_fpAddTest_b_a0_a_a3_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist18_exp_aSig_uid21_fpAddTest_b_2_delay_0_a7_a_aq));
defparam fp_functions_0_aredist18_exp_aSig_uid21_fpAddTest_b_2_delay_0_a7_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist18_exp_aSig_uid21_fpAddTest_b_2_delay_0_a7_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist18_exp_aSig_uid21_fpAddTest_b_2_delay_0_a0_a(
	.clk(clk),
	.d(fp_functions_0_aexp_aSig_uid21_fpAddTest_b_a0_a_a4_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist18_exp_aSig_uid21_fpAddTest_b_2_delay_0_a0_a_aq));
defparam fp_functions_0_aredist18_exp_aSig_uid21_fpAddTest_b_2_delay_0_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist18_exp_aSig_uid21_fpAddTest_b_2_delay_0_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist18_exp_aSig_uid21_fpAddTest_b_2_delay_0_a1_a(
	.clk(clk),
	.d(fp_functions_0_aexp_aSig_uid21_fpAddTest_b_a0_a_a5_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist18_exp_aSig_uid21_fpAddTest_b_2_delay_0_a1_a_aq));
defparam fp_functions_0_aredist18_exp_aSig_uid21_fpAddTest_b_2_delay_0_a1_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist18_exp_aSig_uid21_fpAddTest_b_2_delay_0_a1_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist18_exp_aSig_uid21_fpAddTest_b_2_delay_0_a2_a(
	.clk(clk),
	.d(fp_functions_0_aexp_aSig_uid21_fpAddTest_b_a0_a_a6_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist18_exp_aSig_uid21_fpAddTest_b_2_delay_0_a2_a_aq));
defparam fp_functions_0_aredist18_exp_aSig_uid21_fpAddTest_b_2_delay_0_a2_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist18_exp_aSig_uid21_fpAddTest_b_2_delay_0_a2_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist18_exp_aSig_uid21_fpAddTest_b_2_delay_0_a3_a(
	.clk(clk),
	.d(fp_functions_0_aexp_aSig_uid21_fpAddTest_b_a0_a_a7_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist18_exp_aSig_uid21_fpAddTest_b_2_delay_0_a3_a_aq));
defparam fp_functions_0_aredist18_exp_aSig_uid21_fpAddTest_b_2_delay_0_a3_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist18_exp_aSig_uid21_fpAddTest_b_2_delay_0_a3_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist13_excZ_bSig_uid17_uid37_fpAddTest_q_2_delay_0_a0_a(
	.clk(clk),
	.d(fp_functions_0_areduce_nor_0_a_wirecell_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist13_excZ_bSig_uid17_uid37_fpAddTest_q_2_delay_0_a0_a_aq));
defparam fp_functions_0_aredist13_excZ_bSig_uid17_uid37_fpAddTest_q_2_delay_0_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist13_excZ_bSig_uid17_uid37_fpAddTest_q_2_delay_0_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist7_sigA_uid50_fpAddTest_b_1_q_a0_a(
	.clk(clk),
	.d(fp_functions_0_ai326_a0_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist7_sigA_uid50_fpAddTest_b_1_q_a0_a_aq));
defparam fp_functions_0_aredist7_sigA_uid50_fpAddTest_b_1_q_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist7_sigA_uid50_fpAddTest_b_1_q_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist5_sigB_uid51_fpAddTest_b_1_q_a0_a(
	.clk(clk),
	.d(fp_functions_0_ai289_a0_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist5_sigB_uid51_fpAddTest_b_1_q_a0_a_aq));
defparam fp_functions_0_aredist5_sigB_uid51_fpAddTest_b_1_q_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist5_sigB_uid51_fpAddTest_b_1_q_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist17_frac_aSig_uid22_fpAddTest_b_1_q_a19_a(
	.clk(clk),
	.d(fp_functions_0_ai2131_a0_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist17_frac_aSig_uid22_fpAddTest_b_1_q_a19_a_aq));
defparam fp_functions_0_aredist17_frac_aSig_uid22_fpAddTest_b_1_q_a19_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist17_frac_aSig_uid22_fpAddTest_b_1_q_a19_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist17_frac_aSig_uid22_fpAddTest_b_1_q_a21_a(
	.clk(clk),
	.d(fp_functions_0_ai2131_a1_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist17_frac_aSig_uid22_fpAddTest_b_1_q_a21_a_aq));
defparam fp_functions_0_aredist17_frac_aSig_uid22_fpAddTest_b_1_q_a21_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist17_frac_aSig_uid22_fpAddTest_b_1_q_a21_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist17_frac_aSig_uid22_fpAddTest_b_1_q_a15_a(
	.clk(clk),
	.d(fp_functions_0_ai2131_a2_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist17_frac_aSig_uid22_fpAddTest_b_1_q_a15_a_aq));
defparam fp_functions_0_aredist17_frac_aSig_uid22_fpAddTest_b_1_q_a15_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist17_frac_aSig_uid22_fpAddTest_b_1_q_a15_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist17_frac_aSig_uid22_fpAddTest_b_1_q_a16_a(
	.clk(clk),
	.d(fp_functions_0_ai2131_a3_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist17_frac_aSig_uid22_fpAddTest_b_1_q_a16_a_aq));
defparam fp_functions_0_aredist17_frac_aSig_uid22_fpAddTest_b_1_q_a16_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist17_frac_aSig_uid22_fpAddTest_b_1_q_a16_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist17_frac_aSig_uid22_fpAddTest_b_1_q_a17_a(
	.clk(clk),
	.d(fp_functions_0_ai2131_a4_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist17_frac_aSig_uid22_fpAddTest_b_1_q_a17_a_aq));
defparam fp_functions_0_aredist17_frac_aSig_uid22_fpAddTest_b_1_q_a17_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist17_frac_aSig_uid22_fpAddTest_b_1_q_a17_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist17_frac_aSig_uid22_fpAddTest_b_1_q_a18_a(
	.clk(clk),
	.d(fp_functions_0_ai2131_a5_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist17_frac_aSig_uid22_fpAddTest_b_1_q_a18_a_aq));
defparam fp_functions_0_aredist17_frac_aSig_uid22_fpAddTest_b_1_q_a18_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist17_frac_aSig_uid22_fpAddTest_b_1_q_a18_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist17_frac_aSig_uid22_fpAddTest_b_1_q_a20_a(
	.clk(clk),
	.d(fp_functions_0_ai2131_a6_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist17_frac_aSig_uid22_fpAddTest_b_1_q_a20_a_aq));
defparam fp_functions_0_aredist17_frac_aSig_uid22_fpAddTest_b_1_q_a20_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist17_frac_aSig_uid22_fpAddTest_b_1_q_a20_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist17_frac_aSig_uid22_fpAddTest_b_1_q_a22_a(
	.clk(clk),
	.d(fp_functions_0_ai2131_a7_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist17_frac_aSig_uid22_fpAddTest_b_1_q_a22_a_aq));
defparam fp_functions_0_aredist17_frac_aSig_uid22_fpAddTest_b_1_q_a22_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist17_frac_aSig_uid22_fpAddTest_b_1_q_a22_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist17_frac_aSig_uid22_fpAddTest_b_1_q_a2_a(
	.clk(clk),
	.d(fp_functions_0_ai2131_a8_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist17_frac_aSig_uid22_fpAddTest_b_1_q_a2_a_aq));
defparam fp_functions_0_aredist17_frac_aSig_uid22_fpAddTest_b_1_q_a2_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist17_frac_aSig_uid22_fpAddTest_b_1_q_a2_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist17_frac_aSig_uid22_fpAddTest_b_1_q_a0_a(
	.clk(clk),
	.d(fp_functions_0_ai2131_a9_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist17_frac_aSig_uid22_fpAddTest_b_1_q_a0_a_aq));
defparam fp_functions_0_aredist17_frac_aSig_uid22_fpAddTest_b_1_q_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist17_frac_aSig_uid22_fpAddTest_b_1_q_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist17_frac_aSig_uid22_fpAddTest_b_1_q_a1_a(
	.clk(clk),
	.d(fp_functions_0_ai2131_a10_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist17_frac_aSig_uid22_fpAddTest_b_1_q_a1_a_aq));
defparam fp_functions_0_aredist17_frac_aSig_uid22_fpAddTest_b_1_q_a1_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist17_frac_aSig_uid22_fpAddTest_b_1_q_a1_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist17_frac_aSig_uid22_fpAddTest_b_1_q_a8_a(
	.clk(clk),
	.d(fp_functions_0_ai2131_a11_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist17_frac_aSig_uid22_fpAddTest_b_1_q_a8_a_aq));
defparam fp_functions_0_aredist17_frac_aSig_uid22_fpAddTest_b_1_q_a8_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist17_frac_aSig_uid22_fpAddTest_b_1_q_a8_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist17_frac_aSig_uid22_fpAddTest_b_1_q_a13_a(
	.clk(clk),
	.d(fp_functions_0_ai2131_a12_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist17_frac_aSig_uid22_fpAddTest_b_1_q_a13_a_aq));
defparam fp_functions_0_aredist17_frac_aSig_uid22_fpAddTest_b_1_q_a13_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist17_frac_aSig_uid22_fpAddTest_b_1_q_a13_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist17_frac_aSig_uid22_fpAddTest_b_1_q_a14_a(
	.clk(clk),
	.d(fp_functions_0_ai2131_a13_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist17_frac_aSig_uid22_fpAddTest_b_1_q_a14_a_aq));
defparam fp_functions_0_aredist17_frac_aSig_uid22_fpAddTest_b_1_q_a14_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist17_frac_aSig_uid22_fpAddTest_b_1_q_a14_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist17_frac_aSig_uid22_fpAddTest_b_1_q_a9_a(
	.clk(clk),
	.d(fp_functions_0_ai2131_a14_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist17_frac_aSig_uid22_fpAddTest_b_1_q_a9_a_aq));
defparam fp_functions_0_aredist17_frac_aSig_uid22_fpAddTest_b_1_q_a9_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist17_frac_aSig_uid22_fpAddTest_b_1_q_a9_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist17_frac_aSig_uid22_fpAddTest_b_1_q_a10_a(
	.clk(clk),
	.d(fp_functions_0_ai2131_a15_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist17_frac_aSig_uid22_fpAddTest_b_1_q_a10_a_aq));
defparam fp_functions_0_aredist17_frac_aSig_uid22_fpAddTest_b_1_q_a10_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist17_frac_aSig_uid22_fpAddTest_b_1_q_a10_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist17_frac_aSig_uid22_fpAddTest_b_1_q_a11_a(
	.clk(clk),
	.d(fp_functions_0_ai2131_a16_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist17_frac_aSig_uid22_fpAddTest_b_1_q_a11_a_aq));
defparam fp_functions_0_aredist17_frac_aSig_uid22_fpAddTest_b_1_q_a11_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist17_frac_aSig_uid22_fpAddTest_b_1_q_a11_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist17_frac_aSig_uid22_fpAddTest_b_1_q_a12_a(
	.clk(clk),
	.d(fp_functions_0_ai2131_a17_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist17_frac_aSig_uid22_fpAddTest_b_1_q_a12_a_aq));
defparam fp_functions_0_aredist17_frac_aSig_uid22_fpAddTest_b_1_q_a12_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist17_frac_aSig_uid22_fpAddTest_b_1_q_a12_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist17_frac_aSig_uid22_fpAddTest_b_1_q_a3_a(
	.clk(clk),
	.d(fp_functions_0_ai2131_a18_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist17_frac_aSig_uid22_fpAddTest_b_1_q_a3_a_aq));
defparam fp_functions_0_aredist17_frac_aSig_uid22_fpAddTest_b_1_q_a3_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist17_frac_aSig_uid22_fpAddTest_b_1_q_a3_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist17_frac_aSig_uid22_fpAddTest_b_1_q_a4_a(
	.clk(clk),
	.d(fp_functions_0_ai2131_a19_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist17_frac_aSig_uid22_fpAddTest_b_1_q_a4_a_aq));
defparam fp_functions_0_aredist17_frac_aSig_uid22_fpAddTest_b_1_q_a4_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist17_frac_aSig_uid22_fpAddTest_b_1_q_a4_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist17_frac_aSig_uid22_fpAddTest_b_1_q_a5_a(
	.clk(clk),
	.d(fp_functions_0_ai2131_a20_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist17_frac_aSig_uid22_fpAddTest_b_1_q_a5_a_aq));
defparam fp_functions_0_aredist17_frac_aSig_uid22_fpAddTest_b_1_q_a5_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist17_frac_aSig_uid22_fpAddTest_b_1_q_a5_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist17_frac_aSig_uid22_fpAddTest_b_1_q_a6_a(
	.clk(clk),
	.d(fp_functions_0_ai2131_a21_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist17_frac_aSig_uid22_fpAddTest_b_1_q_a6_a_aq));
defparam fp_functions_0_aredist17_frac_aSig_uid22_fpAddTest_b_1_q_a6_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist17_frac_aSig_uid22_fpAddTest_b_1_q_a6_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist17_frac_aSig_uid22_fpAddTest_b_1_q_a7_a(
	.clk(clk),
	.d(fp_functions_0_ai2131_a22_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist17_frac_aSig_uid22_fpAddTest_b_1_q_a7_a_aq));
defparam fp_functions_0_aredist17_frac_aSig_uid22_fpAddTest_b_1_q_a7_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist17_frac_aSig_uid22_fpAddTest_b_1_q_a7_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_afracXIsZero_uid39_fpAddTest_delay_adelay_signals_a0_a_a0_a(
	.clk(clk),
	.d(fp_functions_0_areduce_nor_10_acombout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_afracXIsZero_uid39_fpAddTest_delay_adelay_signals_a0_a_a0_a_aq));
defparam fp_functions_0_afracXIsZero_uid39_fpAddTest_delay_adelay_signals_a0_a_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_afracXIsZero_uid39_fpAddTest_delay_adelay_signals_a0_a_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist0_vStage_uid154_lzCountVal_uid85_fpAddTest_b_1_q_a0_a(
	.clk(clk),
	.d(fp_functions_0_areduce_nor_1_a4_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist0_vStage_uid154_lzCountVal_uid85_fpAddTest_b_1_q_a0_a_aq));
defparam fp_functions_0_aredist0_vStage_uid154_lzCountVal_uid85_fpAddTest_b_1_q_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist0_vStage_uid154_lzCountVal_uid85_fpAddTest_b_1_q_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist0_vStage_uid154_lzCountVal_uid85_fpAddTest_b_1_q_a3_a(
	.clk(clk),
	.d(fp_functions_0_aadd_4_a111_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist0_vStage_uid154_lzCountVal_uid85_fpAddTest_b_1_q_a3_a_aq));
defparam fp_functions_0_aredist0_vStage_uid154_lzCountVal_uid85_fpAddTest_b_1_q_a3_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist0_vStage_uid154_lzCountVal_uid85_fpAddTest_b_1_q_a3_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist0_vStage_uid154_lzCountVal_uid85_fpAddTest_b_1_q_a1_a(
	.clk(clk),
	.d(fp_functions_0_aadd_4_a131_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist0_vStage_uid154_lzCountVal_uid85_fpAddTest_b_1_q_a1_a_aq));
defparam fp_functions_0_aredist0_vStage_uid154_lzCountVal_uid85_fpAddTest_b_1_q_a1_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist0_vStage_uid154_lzCountVal_uid85_fpAddTest_b_1_q_a1_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist0_vStage_uid154_lzCountVal_uid85_fpAddTest_b_1_q_a4_a(
	.clk(clk),
	.d(fp_functions_0_aadd_4_a91_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist0_vStage_uid154_lzCountVal_uid85_fpAddTest_b_1_q_a4_a_aq));
defparam fp_functions_0_aredist0_vStage_uid154_lzCountVal_uid85_fpAddTest_b_1_q_a4_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist0_vStage_uid154_lzCountVal_uid85_fpAddTest_b_1_q_a4_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist0_vStage_uid154_lzCountVal_uid85_fpAddTest_b_1_q_a2_a(
	.clk(clk),
	.d(fp_functions_0_aadd_4_a126_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist0_vStage_uid154_lzCountVal_uid85_fpAddTest_b_1_q_a2_a_aq));
defparam fp_functions_0_aredist0_vStage_uid154_lzCountVal_uid85_fpAddTest_b_1_q_a2_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist0_vStage_uid154_lzCountVal_uid85_fpAddTest_b_1_q_a2_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aleftShiftStage2_uid249_fracPostNormExt_uid88_fpAddTest_q_a3_a(
	.clk(clk),
	.d(fp_functions_0_ai3337_a3_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aleftShiftStage2_uid249_fracPostNormExt_uid88_fpAddTest_q_a3_a_aq));
defparam fp_functions_0_aleftShiftStage2_uid249_fracPostNormExt_uid88_fpAddTest_q_a3_a.is_wysiwyg = "true";
defparam fp_functions_0_aleftShiftStage2_uid249_fracPostNormExt_uid88_fpAddTest_q_a3_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aleftShiftStage2_uid249_fracPostNormExt_uid88_fpAddTest_q_a2_a(
	.clk(clk),
	.d(fp_functions_0_ai3337_a5_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aleftShiftStage2_uid249_fracPostNormExt_uid88_fpAddTest_q_a2_a_aq));
defparam fp_functions_0_aleftShiftStage2_uid249_fracPostNormExt_uid88_fpAddTest_q_a2_a.is_wysiwyg = "true";
defparam fp_functions_0_aleftShiftStage2_uid249_fracPostNormExt_uid88_fpAddTest_q_a2_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aleftShiftStage2_uid249_fracPostNormExt_uid88_fpAddTest_q_a0_a(
	.clk(clk),
	.d(fp_functions_0_ai3337_a6_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aleftShiftStage2_uid249_fracPostNormExt_uid88_fpAddTest_q_a0_a_aq));
defparam fp_functions_0_aleftShiftStage2_uid249_fracPostNormExt_uid88_fpAddTest_q_a0_a.is_wysiwyg = "true";
defparam fp_functions_0_aleftShiftStage2_uid249_fracPostNormExt_uid88_fpAddTest_q_a0_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aleftShiftStage2_uid249_fracPostNormExt_uid88_fpAddTest_q_a1_a(
	.clk(clk),
	.d(fp_functions_0_ai3337_a7_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aleftShiftStage2_uid249_fracPostNormExt_uid88_fpAddTest_q_a1_a_aq));
defparam fp_functions_0_aleftShiftStage2_uid249_fracPostNormExt_uid88_fpAddTest_q_a1_a.is_wysiwyg = "true";
defparam fp_functions_0_aleftShiftStage2_uid249_fracPostNormExt_uid88_fpAddTest_q_a1_a.power_up = "dont_care";

fourteennm_lcell_comb fp_functions_0_aadd_6_a1(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!fp_functions_0_aadd_5_a1_sumout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_6_a27),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_6_a1_sumout),
	.cout(fp_functions_0_aadd_6_a2),
	.shareout());
defparam fp_functions_0_aadd_6_a1.extended_lut = "off";
defparam fp_functions_0_aadd_6_a1.lut_mask = 64'h0000000000FFFF00;
defparam fp_functions_0_aadd_6_a1.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_6_a6(
	.dataa(!fp_functions_0_arVStage_uid165_lzCountVal_uid85_fpAddTest_merged_bit_select_b_a3_a_a6_combout),
	.datab(!fp_functions_0_arVStage_uid177_lzCountVal_uid85_fpAddTest_b_a0_a_a0_combout),
	.datac(!fp_functions_0_arVStage_uid171_lzCountVal_uid85_fpAddTest_merged_bit_select_b_a1_a_a3_combout),
	.datad(!fp_functions_0_aadd_5_a6_sumout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_6_a52_cout),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_6_a6_sumout),
	.cout(fp_functions_0_aadd_6_a7),
	.shareout());
defparam fp_functions_0_aadd_6_a6.extended_lut = "off";
defparam fp_functions_0_aadd_6_a6.lut_mask = 64'h0000000000BFBF40;
defparam fp_functions_0_aadd_6_a6.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_6_a11(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_areduce_nor_5_a0_combout),
	.datad(!fp_functions_0_aadd_5_a11_sumout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_6_a7),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_6_a11_sumout),
	.cout(fp_functions_0_aadd_6_a12),
	.shareout());
defparam fp_functions_0_aadd_6_a11.extended_lut = "off";
defparam fp_functions_0_aadd_6_a11.lut_mask = 64'h00000000000F0FF0;
defparam fp_functions_0_aadd_6_a11.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_6_a16(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_areduce_nor_4_acombout),
	.datad(!fp_functions_0_aadd_5_a16_sumout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_6_a12),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_6_a16_sumout),
	.cout(fp_functions_0_aadd_6_a17),
	.shareout());
defparam fp_functions_0_aadd_6_a16.extended_lut = "off";
defparam fp_functions_0_aadd_6_a16.lut_mask = 64'h00000000000F0FF0;
defparam fp_functions_0_aadd_6_a16.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_6_a21(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_areduce_nor_3_acombout),
	.datad(!fp_functions_0_aadd_5_a21_sumout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_6_a17),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_6_a21_sumout),
	.cout(fp_functions_0_aadd_6_a22),
	.shareout());
defparam fp_functions_0_aadd_6_a21.extended_lut = "off";
defparam fp_functions_0_aadd_6_a21.lut_mask = 64'h00000000000F0FF0;
defparam fp_functions_0_aadd_6_a21.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_6_a26(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aredist1_vCount_uid152_lzCountVal_uid85_fpAddTest_q_1_q_a0_a_aq),
	.datad(!fp_functions_0_aadd_5_a26_sumout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_6_a22),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_6_a26_sumout),
	.cout(fp_functions_0_aadd_6_a27),
	.shareout());
defparam fp_functions_0_aadd_6_a26.extended_lut = "off";
defparam fp_functions_0_aadd_6_a26.lut_mask = 64'h0000000000F0F00F;
defparam fp_functions_0_aadd_6_a26.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_6_a31(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!fp_functions_0_aadd_5_a31_sumout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_6_a2),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_6_a31_sumout),
	.cout(fp_functions_0_aadd_6_a32),
	.shareout());
defparam fp_functions_0_aadd_6_a31.extended_lut = "off";
defparam fp_functions_0_aadd_6_a31.lut_mask = 64'h0000000000FFFF00;
defparam fp_functions_0_aadd_6_a31.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_6_a36(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!fp_functions_0_aadd_5_a36_sumout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_6_a32),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_6_a36_sumout),
	.cout(fp_functions_0_aadd_6_a37),
	.shareout());
defparam fp_functions_0_aadd_6_a36.extended_lut = "off";
defparam fp_functions_0_aadd_6_a36.lut_mask = 64'h0000000000FFFF00;
defparam fp_functions_0_aadd_6_a36.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_6_a41(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!fp_functions_0_aadd_5_a41_sumout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_6_a37),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_6_a41_sumout),
	.cout(fp_functions_0_aadd_6_a42),
	.shareout());
defparam fp_functions_0_aadd_6_a41.extended_lut = "off";
defparam fp_functions_0_aadd_6_a41.lut_mask = 64'h0000000000FFFF00;
defparam fp_functions_0_aadd_6_a41.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_6_a46(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_6_a42),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_6_a46_sumout),
	.cout(),
	.shareout());
defparam fp_functions_0_aadd_6_a46.extended_lut = "off";
defparam fp_functions_0_aadd_6_a46.lut_mask = 64'h000000000000FFFF;
defparam fp_functions_0_aadd_6_a46.shared_arith = "off";

fourteennm_ff fp_functions_0_aredist0_vStage_uid154_lzCountVal_uid85_fpAddTest_b_1_q_a5_a(
	.clk(clk),
	.d(fp_functions_0_aadd_4_a96_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist0_vStage_uid154_lzCountVal_uid85_fpAddTest_b_1_q_a5_a_aq));
defparam fp_functions_0_aredist0_vStage_uid154_lzCountVal_uid85_fpAddTest_b_1_q_a5_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist0_vStage_uid154_lzCountVal_uid85_fpAddTest_b_1_q_a5_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist0_vStage_uid154_lzCountVal_uid85_fpAddTest_b_1_q_a6_a(
	.clk(clk),
	.d(fp_functions_0_aadd_4_a86_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist0_vStage_uid154_lzCountVal_uid85_fpAddTest_b_1_q_a6_a_aq));
defparam fp_functions_0_aredist0_vStage_uid154_lzCountVal_uid85_fpAddTest_b_1_q_a6_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist0_vStage_uid154_lzCountVal_uid85_fpAddTest_b_1_q_a6_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist0_vStage_uid154_lzCountVal_uid85_fpAddTest_b_1_q_a7_a(
	.clk(clk),
	.d(fp_functions_0_aadd_4_a81_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist0_vStage_uid154_lzCountVal_uid85_fpAddTest_b_1_q_a7_a_aq));
defparam fp_functions_0_aredist0_vStage_uid154_lzCountVal_uid85_fpAddTest_b_1_q_a7_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist0_vStage_uid154_lzCountVal_uid85_fpAddTest_b_1_q_a7_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist0_vStage_uid154_lzCountVal_uid85_fpAddTest_b_1_q_a8_a(
	.clk(clk),
	.d(fp_functions_0_aadd_4_a116_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist0_vStage_uid154_lzCountVal_uid85_fpAddTest_b_1_q_a8_a_aq));
defparam fp_functions_0_aredist0_vStage_uid154_lzCountVal_uid85_fpAddTest_b_1_q_a8_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist0_vStage_uid154_lzCountVal_uid85_fpAddTest_b_1_q_a8_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist0_vStage_uid154_lzCountVal_uid85_fpAddTest_b_1_q_a9_a(
	.clk(clk),
	.d(fp_functions_0_aadd_4_a121_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist0_vStage_uid154_lzCountVal_uid85_fpAddTest_b_1_q_a9_a_aq));
defparam fp_functions_0_aredist0_vStage_uid154_lzCountVal_uid85_fpAddTest_b_1_q_a9_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist0_vStage_uid154_lzCountVal_uid85_fpAddTest_b_1_q_a9_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist0_vStage_uid154_lzCountVal_uid85_fpAddTest_b_1_q_a10_a(
	.clk(clk),
	.d(fp_functions_0_aadd_4_a106_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist0_vStage_uid154_lzCountVal_uid85_fpAddTest_b_1_q_a10_a_aq));
defparam fp_functions_0_aredist0_vStage_uid154_lzCountVal_uid85_fpAddTest_b_1_q_a10_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist0_vStage_uid154_lzCountVal_uid85_fpAddTest_b_1_q_a10_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist3_fracGRS_uid84_fpAddTest_q_1_q_a11_a(
	.clk(clk),
	.d(fp_functions_0_aadd_4_a101_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist3_fracGRS_uid84_fpAddTest_q_1_q_a11_a_aq));
defparam fp_functions_0_aredist3_fracGRS_uid84_fpAddTest_q_1_q_a11_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist3_fracGRS_uid84_fpAddTest_q_1_q_a11_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist3_fracGRS_uid84_fpAddTest_q_1_q_a12_a(
	.clk(clk),
	.d(fp_functions_0_aadd_4_a11_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist3_fracGRS_uid84_fpAddTest_q_1_q_a12_a_aq));
defparam fp_functions_0_aredist3_fracGRS_uid84_fpAddTest_q_1_q_a12_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist3_fracGRS_uid84_fpAddTest_q_1_q_a12_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist3_fracGRS_uid84_fpAddTest_q_1_q_a13_a(
	.clk(clk),
	.d(fp_functions_0_aadd_4_a16_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist3_fracGRS_uid84_fpAddTest_q_1_q_a13_a_aq));
defparam fp_functions_0_aredist3_fracGRS_uid84_fpAddTest_q_1_q_a13_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist3_fracGRS_uid84_fpAddTest_q_1_q_a13_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist3_fracGRS_uid84_fpAddTest_q_1_q_a14_a(
	.clk(clk),
	.d(fp_functions_0_aadd_4_a21_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist3_fracGRS_uid84_fpAddTest_q_1_q_a14_a_aq));
defparam fp_functions_0_aredist3_fracGRS_uid84_fpAddTest_q_1_q_a14_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist3_fracGRS_uid84_fpAddTest_q_1_q_a14_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist3_fracGRS_uid84_fpAddTest_q_1_q_a15_a(
	.clk(clk),
	.d(fp_functions_0_aadd_4_a26_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist3_fracGRS_uid84_fpAddTest_q_1_q_a15_a_aq));
defparam fp_functions_0_aredist3_fracGRS_uid84_fpAddTest_q_1_q_a15_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist3_fracGRS_uid84_fpAddTest_q_1_q_a15_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist3_fracGRS_uid84_fpAddTest_q_1_q_a16_a(
	.clk(clk),
	.d(fp_functions_0_aadd_4_a6_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist3_fracGRS_uid84_fpAddTest_q_1_q_a16_a_aq));
defparam fp_functions_0_aredist3_fracGRS_uid84_fpAddTest_q_1_q_a16_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist3_fracGRS_uid84_fpAddTest_q_1_q_a16_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist3_fracGRS_uid84_fpAddTest_q_1_q_a17_a(
	.clk(clk),
	.d(fp_functions_0_aadd_4_a31_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist3_fracGRS_uid84_fpAddTest_q_1_q_a17_a_aq));
defparam fp_functions_0_aredist3_fracGRS_uid84_fpAddTest_q_1_q_a17_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist3_fracGRS_uid84_fpAddTest_q_1_q_a17_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist3_fracGRS_uid84_fpAddTest_q_1_q_a18_a(
	.clk(clk),
	.d(fp_functions_0_aadd_4_a36_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist3_fracGRS_uid84_fpAddTest_q_1_q_a18_a_aq));
defparam fp_functions_0_aredist3_fracGRS_uid84_fpAddTest_q_1_q_a18_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist3_fracGRS_uid84_fpAddTest_q_1_q_a18_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist3_fracGRS_uid84_fpAddTest_q_1_q_a19_a(
	.clk(clk),
	.d(fp_functions_0_aadd_4_a41_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist3_fracGRS_uid84_fpAddTest_q_1_q_a19_a_aq));
defparam fp_functions_0_aredist3_fracGRS_uid84_fpAddTest_q_1_q_a19_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist3_fracGRS_uid84_fpAddTest_q_1_q_a19_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist3_fracGRS_uid84_fpAddTest_q_1_q_a20_a(
	.clk(clk),
	.d(fp_functions_0_aadd_4_a1_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist3_fracGRS_uid84_fpAddTest_q_1_q_a20_a_aq));
defparam fp_functions_0_aredist3_fracGRS_uid84_fpAddTest_q_1_q_a20_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist3_fracGRS_uid84_fpAddTest_q_1_q_a20_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist3_fracGRS_uid84_fpAddTest_q_1_q_a21_a(
	.clk(clk),
	.d(fp_functions_0_aadd_4_a56_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist3_fracGRS_uid84_fpAddTest_q_1_q_a21_a_aq));
defparam fp_functions_0_aredist3_fracGRS_uid84_fpAddTest_q_1_q_a21_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist3_fracGRS_uid84_fpAddTest_q_1_q_a21_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist3_fracGRS_uid84_fpAddTest_q_1_q_a22_a(
	.clk(clk),
	.d(fp_functions_0_aadd_4_a61_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist3_fracGRS_uid84_fpAddTest_q_1_q_a22_a_aq));
defparam fp_functions_0_aredist3_fracGRS_uid84_fpAddTest_q_1_q_a22_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist3_fracGRS_uid84_fpAddTest_q_1_q_a22_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist3_fracGRS_uid84_fpAddTest_q_1_q_a23_a(
	.clk(clk),
	.d(fp_functions_0_aadd_4_a66_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist3_fracGRS_uid84_fpAddTest_q_1_q_a23_a_aq));
defparam fp_functions_0_aredist3_fracGRS_uid84_fpAddTest_q_1_q_a23_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist3_fracGRS_uid84_fpAddTest_q_1_q_a23_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist3_fracGRS_uid84_fpAddTest_q_1_q_a24_a(
	.clk(clk),
	.d(fp_functions_0_aadd_4_a71_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist3_fracGRS_uid84_fpAddTest_q_1_q_a24_a_aq));
defparam fp_functions_0_aredist3_fracGRS_uid84_fpAddTest_q_1_q_a24_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist3_fracGRS_uid84_fpAddTest_q_1_q_a24_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist3_fracGRS_uid84_fpAddTest_q_1_q_a25_a(
	.clk(clk),
	.d(fp_functions_0_aadd_4_a46_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist3_fracGRS_uid84_fpAddTest_q_1_q_a25_a_aq));
defparam fp_functions_0_aredist3_fracGRS_uid84_fpAddTest_q_1_q_a25_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist3_fracGRS_uid84_fpAddTest_q_1_q_a25_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_aredist3_fracGRS_uid84_fpAddTest_q_1_q_a26_a(
	.clk(clk),
	.d(fp_functions_0_aadd_4_a51_sumout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(areset),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_aredist3_fracGRS_uid84_fpAddTest_q_1_q_a26_a_aq));
defparam fp_functions_0_aredist3_fracGRS_uid84_fpAddTest_q_1_q_a26_a.is_wysiwyg = "true";
defparam fp_functions_0_aredist3_fracGRS_uid84_fpAddTest_q_1_q_a26_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a42_a(
	.clk(clk),
	.d(fp_functions_0_aMux_55_a1_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a41_a_a3_combout),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a42_a_aq));
defparam fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a42_a.is_wysiwyg = "true";
defparam fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a42_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a38_a(
	.clk(clk),
	.d(fp_functions_0_aMux_59_a7_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a41_a_a3_combout),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a38_a_aq));
defparam fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a38_a.is_wysiwyg = "true";
defparam fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a38_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a34_a(
	.clk(clk),
	.d(fp_functions_0_aMux_63_a0_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a41_a_a3_combout),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a34_a_aq));
defparam fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a34_a.is_wysiwyg = "true";
defparam fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a34_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a35_a(
	.clk(clk),
	.d(fp_functions_0_aMux_62_a1_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a41_a_a3_combout),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a35_a_aq));
defparam fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a35_a.is_wysiwyg = "true";
defparam fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a35_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a36_a(
	.clk(clk),
	.d(fp_functions_0_aMux_61_a1_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a41_a_a3_combout),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a36_a_aq));
defparam fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a36_a.is_wysiwyg = "true";
defparam fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a36_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a37_a(
	.clk(clk),
	.d(fp_functions_0_aMux_60_a6_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a41_a_a3_combout),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a37_a_aq));
defparam fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a37_a.is_wysiwyg = "true";
defparam fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a37_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a39_a(
	.clk(clk),
	.d(fp_functions_0_aMux_58_a5_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a41_a_a3_combout),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a39_a_aq));
defparam fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a39_a.is_wysiwyg = "true";
defparam fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a39_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a40_a(
	.clk(clk),
	.d(fp_functions_0_aMux_57_a6_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a41_a_a3_combout),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a40_a_aq));
defparam fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a40_a.is_wysiwyg = "true";
defparam fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a40_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a41_a(
	.clk(clk),
	.d(fp_functions_0_aMux_56_a1_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a41_a_a3_combout),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a41_a_aq));
defparam fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a41_a.is_wysiwyg = "true";
defparam fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a41_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a47_a(
	.clk(clk),
	.d(fp_functions_0_aMux_50_a0_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a41_a_a3_combout),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a47_a_aq));
defparam fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a47_a.is_wysiwyg = "true";
defparam fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a47_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a48_a(
	.clk(clk),
	.d(fp_functions_0_aMux_49_a0_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a41_a_a3_combout),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a48_a_aq));
defparam fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a48_a.is_wysiwyg = "true";
defparam fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a48_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a43_a(
	.clk(clk),
	.d(fp_functions_0_aMux_54_a1_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a41_a_a3_combout),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a43_a_aq));
defparam fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a43_a.is_wysiwyg = "true";
defparam fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a43_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a44_a(
	.clk(clk),
	.d(fp_functions_0_aMux_53_a1_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a41_a_a3_combout),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a44_a_aq));
defparam fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a44_a.is_wysiwyg = "true";
defparam fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a44_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a45_a(
	.clk(clk),
	.d(fp_functions_0_aMux_52_a0_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a41_a_a3_combout),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a45_a_aq));
defparam fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a45_a.is_wysiwyg = "true";
defparam fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a45_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a46_a(
	.clk(clk),
	.d(fp_functions_0_aMux_51_a0_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a41_a_a3_combout),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a46_a_aq));
defparam fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a46_a.is_wysiwyg = "true";
defparam fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a46_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a29_a(
	.clk(clk),
	.d(fp_functions_0_ai1783_a20_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a28_a_a0_combout),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a29_a_aq));
defparam fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a29_a.is_wysiwyg = "true";
defparam fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a29_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a28_a(
	.clk(clk),
	.d(fp_functions_0_ai1783_a21_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a28_a_a0_combout),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a28_a_aq));
defparam fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a28_a.is_wysiwyg = "true";
defparam fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a28_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a26_a(
	.clk(clk),
	.d(fp_functions_0_ai1783_a22_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a28_a_a0_combout),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a26_a_aq));
defparam fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a26_a.is_wysiwyg = "true";
defparam fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a26_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a27_a(
	.clk(clk),
	.d(fp_functions_0_ai1783_a23_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a28_a_a0_combout),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a27_a_aq));
defparam fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a27_a.is_wysiwyg = "true";
defparam fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a27_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a33_a(
	.clk(clk),
	.d(fp_functions_0_aMux_64_a0_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a41_a_a3_combout),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a33_a_aq));
defparam fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a33_a.is_wysiwyg = "true";
defparam fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a33_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a32_a(
	.clk(clk),
	.d(fp_functions_0_ai1783_a24_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a28_a_a0_combout),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a32_a_aq));
defparam fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a32_a.is_wysiwyg = "true";
defparam fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a32_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a25_a(
	.clk(clk),
	.d(fp_functions_0_ai1783_a25_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a28_a_a0_combout),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a25_a_aq));
defparam fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a25_a.is_wysiwyg = "true";
defparam fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a25_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a30_a(
	.clk(clk),
	.d(fp_functions_0_ai1783_a26_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a28_a_a0_combout),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a30_a_aq));
defparam fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a30_a.is_wysiwyg = "true";
defparam fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a30_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a31_a(
	.clk(clk),
	.d(fp_functions_0_ai1783_a27_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a28_a_a0_combout),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a31_a_aq));
defparam fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a31_a.is_wysiwyg = "true";
defparam fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a31_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a24_a(
	.clk(clk),
	.d(fp_functions_0_ai1783_a28_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a28_a_a0_combout),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a24_a_aq));
defparam fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a24_a.is_wysiwyg = "true";
defparam fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a24_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a23_a(
	.clk(clk),
	.d(fp_functions_0_ai1783_a29_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a28_a_a0_combout),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a23_a_aq));
defparam fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a23_a.is_wysiwyg = "true";
defparam fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a23_a.power_up = "dont_care";

fourteennm_lcell_comb fp_functions_0_aadd_2_a1(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_2_a7_cout),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_2_a1_sumout),
	.cout(),
	.shareout());
defparam fp_functions_0_aadd_2_a1.extended_lut = "off";
defparam fp_functions_0_aadd_2_a1.lut_mask = 64'h000000000000FFFF;
defparam fp_functions_0_aadd_2_a1.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_1_a1(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aexp_bSig_uid35_fpAddTest_b_a3_a_a0_combout),
	.datad(!fp_functions_0_aexp_aSig_uid21_fpAddTest_b_a0_a_a7_combout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_1_a22),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_1_a1_sumout),
	.cout(fp_functions_0_aadd_1_a2),
	.shareout());
defparam fp_functions_0_aadd_1_a1.extended_lut = "off";
defparam fp_functions_0_aadd_1_a1.lut_mask = 64'h0000000000F0F00F;
defparam fp_functions_0_aadd_1_a1.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_1_a6(
	.dataa(!fp_functions_0_aadd_0_a1_sumout),
	.datab(!b[27]),
	.datac(!a[27]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_1_a2),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_1_a6_sumout),
	.cout(fp_functions_0_aadd_1_a7),
	.shareout());
defparam fp_functions_0_aadd_1_a6.extended_lut = "off";
defparam fp_functions_0_aadd_1_a6.lut_mask = 64'h000000001818C3C3;
defparam fp_functions_0_aadd_1_a6.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_1_a11(
	.dataa(!fp_functions_0_aadd_0_a1_sumout),
	.datab(!b[23]),
	.datac(!a[23]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_1_a32_cout),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_1_a11_sumout),
	.cout(fp_functions_0_aadd_1_a12),
	.shareout());
defparam fp_functions_0_aadd_1_a11.extended_lut = "off";
defparam fp_functions_0_aadd_1_a11.lut_mask = 64'h000000001818C3C3;
defparam fp_functions_0_aadd_1_a11.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_0_a1(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_0_a7_cout),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_0_a1_sumout),
	.cout(),
	.shareout());
defparam fp_functions_0_aadd_0_a1.extended_lut = "off";
defparam fp_functions_0_aadd_0_a1.lut_mask = 64'h000000000000FFFF;
defparam fp_functions_0_aadd_0_a1.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_1_a16(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aexp_bSig_uid35_fpAddTest_b_a1_a_a1_combout),
	.datad(!fp_functions_0_aexp_aSig_uid21_fpAddTest_b_a0_a_a5_combout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_1_a12),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_1_a16_sumout),
	.cout(fp_functions_0_aadd_1_a17),
	.shareout());
defparam fp_functions_0_aadd_1_a16.extended_lut = "off";
defparam fp_functions_0_aadd_1_a16.lut_mask = 64'h0000000000F0F00F;
defparam fp_functions_0_aadd_1_a16.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_1_a21(
	.dataa(!fp_functions_0_aadd_0_a1_sumout),
	.datab(!b[25]),
	.datac(!a[25]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_1_a17),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_1_a21_sumout),
	.cout(fp_functions_0_aadd_1_a22),
	.shareout());
defparam fp_functions_0_aadd_1_a21.extended_lut = "off";
defparam fp_functions_0_aadd_1_a21.lut_mask = 64'h000000001818C3C3;
defparam fp_functions_0_aadd_1_a21.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_1_a26(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aexp_bSig_uid35_fpAddTest_b_a5_a_a2_combout),
	.datad(!fp_functions_0_aexp_aSig_uid21_fpAddTest_b_a0_a_a1_combout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_1_a7),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_1_a26_sumout),
	.cout(fp_functions_0_aadd_1_a27),
	.shareout());
defparam fp_functions_0_aadd_1_a26.extended_lut = "off";
defparam fp_functions_0_aadd_1_a26.lut_mask = 64'h0000000000F0F00F;
defparam fp_functions_0_aadd_1_a26.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_3_a1(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_3_a7_cout),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_3_a1_sumout),
	.cout(),
	.shareout());
defparam fp_functions_0_aadd_3_a1.extended_lut = "off";
defparam fp_functions_0_aadd_3_a1.lut_mask = 64'h000000000000FFFF;
defparam fp_functions_0_aadd_3_a1.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_5_a1(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aredist18_exp_aSig_uid21_fpAddTest_b_2_q_a5_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_5_a27),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_5_a1_sumout),
	.cout(fp_functions_0_aadd_5_a2),
	.shareout());
defparam fp_functions_0_aadd_5_a1.extended_lut = "off";
defparam fp_functions_0_aadd_5_a1.lut_mask = 64'h0000000000000F0F;
defparam fp_functions_0_aadd_5_a1.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_5_a6(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aredist18_exp_aSig_uid21_fpAddTest_b_2_q_a0_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_5_a6_sumout),
	.cout(fp_functions_0_aadd_5_a7),
	.shareout());
defparam fp_functions_0_aadd_5_a6.extended_lut = "off";
defparam fp_functions_0_aadd_5_a6.lut_mask = 64'h000000000F0FF0F0;
defparam fp_functions_0_aadd_5_a6.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_6_a52(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fp_functions_0_aadd_6_a52_cout),
	.shareout());
defparam fp_functions_0_aadd_6_a52.extended_lut = "off";
defparam fp_functions_0_aadd_6_a52.lut_mask = 64'h00000000FFFF0000;
defparam fp_functions_0_aadd_6_a52.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_5_a11(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aredist18_exp_aSig_uid21_fpAddTest_b_2_q_a1_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_5_a7),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_5_a11_sumout),
	.cout(fp_functions_0_aadd_5_a12),
	.shareout());
defparam fp_functions_0_aadd_5_a11.extended_lut = "off";
defparam fp_functions_0_aadd_5_a11.lut_mask = 64'h0000000000000F0F;
defparam fp_functions_0_aadd_5_a11.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_5_a16(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aredist18_exp_aSig_uid21_fpAddTest_b_2_q_a2_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_5_a12),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_5_a16_sumout),
	.cout(fp_functions_0_aadd_5_a17),
	.shareout());
defparam fp_functions_0_aadd_5_a16.extended_lut = "off";
defparam fp_functions_0_aadd_5_a16.lut_mask = 64'h0000000000000F0F;
defparam fp_functions_0_aadd_5_a16.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_5_a21(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aredist18_exp_aSig_uid21_fpAddTest_b_2_q_a3_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_5_a17),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_5_a21_sumout),
	.cout(fp_functions_0_aadd_5_a22),
	.shareout());
defparam fp_functions_0_aadd_5_a21.extended_lut = "off";
defparam fp_functions_0_aadd_5_a21.lut_mask = 64'h0000000000000F0F;
defparam fp_functions_0_aadd_5_a21.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_5_a26(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aredist18_exp_aSig_uid21_fpAddTest_b_2_q_a4_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_5_a22),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_5_a26_sumout),
	.cout(fp_functions_0_aadd_5_a27),
	.shareout());
defparam fp_functions_0_aadd_5_a26.extended_lut = "off";
defparam fp_functions_0_aadd_5_a26.lut_mask = 64'h0000000000000F0F;
defparam fp_functions_0_aadd_5_a26.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_5_a31(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aredist18_exp_aSig_uid21_fpAddTest_b_2_q_a6_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_5_a2),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_5_a31_sumout),
	.cout(fp_functions_0_aadd_5_a32),
	.shareout());
defparam fp_functions_0_aadd_5_a31.extended_lut = "off";
defparam fp_functions_0_aadd_5_a31.lut_mask = 64'h0000000000000F0F;
defparam fp_functions_0_aadd_5_a31.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_5_a36(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aredist18_exp_aSig_uid21_fpAddTest_b_2_q_a7_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_5_a32),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_5_a36_sumout),
	.cout(fp_functions_0_aadd_5_a37),
	.shareout());
defparam fp_functions_0_aadd_5_a36.extended_lut = "off";
defparam fp_functions_0_aadd_5_a36.lut_mask = 64'h0000000000000F0F;
defparam fp_functions_0_aadd_5_a36.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_5_a41(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_5_a37),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_5_a41_sumout),
	.cout(),
	.shareout());
defparam fp_functions_0_aadd_5_a41.extended_lut = "off";
defparam fp_functions_0_aadd_5_a41.lut_mask = 64'h0000000000000000;
defparam fp_functions_0_aadd_5_a41.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_2_a7(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aadd_1_a36_sumout),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_2_a12_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fp_functions_0_aadd_2_a7_cout),
	.shareout());
defparam fp_functions_0_aadd_2_a7.extended_lut = "off";
defparam fp_functions_0_aadd_2_a7.lut_mask = 64'h000000000000F0F0;
defparam fp_functions_0_aadd_2_a7.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_1_a32(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fp_functions_0_aadd_1_a32_cout),
	.shareout());
defparam fp_functions_0_aadd_1_a32.extended_lut = "off";
defparam fp_functions_0_aadd_1_a32.lut_mask = 64'h00000000FFFF0000;
defparam fp_functions_0_aadd_1_a32.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_0_a7(
	.dataa(gnd),
	.datab(gnd),
	.datac(!b[30]),
	.datad(!a[30]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_0_a12_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fp_functions_0_aadd_0_a7_cout),
	.shareout());
defparam fp_functions_0_aadd_0_a7.extended_lut = "off";
defparam fp_functions_0_aadd_0_a7.lut_mask = 64'h0000000000F0F00F;
defparam fp_functions_0_aadd_0_a7.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_3_a7(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aadd_1_a36_sumout),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_3_a12_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fp_functions_0_aadd_3_a7_cout),
	.shareout());
defparam fp_functions_0_aadd_3_a7.extended_lut = "off";
defparam fp_functions_0_aadd_3_a7.lut_mask = 64'h000000000F0FF0F0;
defparam fp_functions_0_aadd_3_a7.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_1_a36(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_1_a42),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_1_a36_sumout),
	.cout(),
	.shareout());
defparam fp_functions_0_aadd_1_a36.extended_lut = "off";
defparam fp_functions_0_aadd_1_a36.lut_mask = 64'h000000000000FFFF;
defparam fp_functions_0_aadd_1_a36.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_2_a12(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aadd_1_a41_sumout),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_2_a17_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fp_functions_0_aadd_2_a12_cout),
	.shareout());
defparam fp_functions_0_aadd_2_a12.extended_lut = "off";
defparam fp_functions_0_aadd_2_a12.lut_mask = 64'h000000000000F0F0;
defparam fp_functions_0_aadd_2_a12.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_0_a12(
	.dataa(gnd),
	.datab(gnd),
	.datac(!b[29]),
	.datad(!a[29]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_0_a17_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fp_functions_0_aadd_0_a12_cout),
	.shareout());
defparam fp_functions_0_aadd_0_a12.extended_lut = "off";
defparam fp_functions_0_aadd_0_a12.lut_mask = 64'h0000000000F0F00F;
defparam fp_functions_0_aadd_0_a12.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_3_a12(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aadd_1_a41_sumout),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_3_a17_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fp_functions_0_aadd_3_a12_cout),
	.shareout());
defparam fp_functions_0_aadd_3_a12.extended_lut = "off";
defparam fp_functions_0_aadd_3_a12.lut_mask = 64'h000000000F0FF0F0;
defparam fp_functions_0_aadd_3_a12.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_1_a41(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aexp_bSig_uid35_fpAddTest_b_a7_a_a3_combout),
	.datad(!fp_functions_0_aexp_aSig_uid21_fpAddTest_b_a0_a_a3_combout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_1_a47),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_1_a41_sumout),
	.cout(fp_functions_0_aadd_1_a42),
	.shareout());
defparam fp_functions_0_aadd_1_a41.extended_lut = "off";
defparam fp_functions_0_aadd_1_a41.lut_mask = 64'h0000000000F0F00F;
defparam fp_functions_0_aadd_1_a41.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_2_a17(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aadd_1_a46_sumout),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_2_a22_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fp_functions_0_aadd_2_a17_cout),
	.shareout());
defparam fp_functions_0_aadd_2_a17.extended_lut = "off";
defparam fp_functions_0_aadd_2_a17.lut_mask = 64'h000000000000F0F0;
defparam fp_functions_0_aadd_2_a17.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_0_a17(
	.dataa(gnd),
	.datab(gnd),
	.datac(!b[28]),
	.datad(!a[28]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_0_a22_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fp_functions_0_aadd_0_a17_cout),
	.shareout());
defparam fp_functions_0_aadd_0_a17.extended_lut = "off";
defparam fp_functions_0_aadd_0_a17.lut_mask = 64'h0000000000F0F00F;
defparam fp_functions_0_aadd_0_a17.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_3_a17(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aadd_1_a46_sumout),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_3_a22_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fp_functions_0_aadd_3_a17_cout),
	.shareout());
defparam fp_functions_0_aadd_3_a17.extended_lut = "off";
defparam fp_functions_0_aadd_3_a17.lut_mask = 64'h000000000F0FF0F0;
defparam fp_functions_0_aadd_3_a17.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_1_a46(
	.dataa(!fp_functions_0_aadd_0_a1_sumout),
	.datab(!b[29]),
	.datac(!a[29]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_1_a27),
	.sharein(gnd),
	.combout(),
	.sumout(fp_functions_0_aadd_1_a46_sumout),
	.cout(fp_functions_0_aadd_1_a47),
	.shareout());
defparam fp_functions_0_aadd_1_a46.extended_lut = "off";
defparam fp_functions_0_aadd_1_a46.lut_mask = 64'h000000001818C3C3;
defparam fp_functions_0_aadd_1_a46.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_2_a22(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aadd_1_a26_sumout),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_2_a27_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fp_functions_0_aadd_2_a22_cout),
	.shareout());
defparam fp_functions_0_aadd_2_a22.extended_lut = "off";
defparam fp_functions_0_aadd_2_a22.lut_mask = 64'h000000000000F0F0;
defparam fp_functions_0_aadd_2_a22.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_0_a22(
	.dataa(gnd),
	.datab(gnd),
	.datac(!b[27]),
	.datad(!a[27]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_0_a27_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fp_functions_0_aadd_0_a22_cout),
	.shareout());
defparam fp_functions_0_aadd_0_a22.extended_lut = "off";
defparam fp_functions_0_aadd_0_a22.lut_mask = 64'h0000000000F0F00F;
defparam fp_functions_0_aadd_0_a22.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_3_a22(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aadd_1_a26_sumout),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_3_a27_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fp_functions_0_aadd_3_a22_cout),
	.shareout());
defparam fp_functions_0_aadd_3_a22.extended_lut = "off";
defparam fp_functions_0_aadd_3_a22.lut_mask = 64'h0000000000000F0F;
defparam fp_functions_0_aadd_3_a22.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_2_a27(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aadd_1_a6_sumout),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_2_a32_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fp_functions_0_aadd_2_a27_cout),
	.shareout());
defparam fp_functions_0_aadd_2_a27.extended_lut = "off";
defparam fp_functions_0_aadd_2_a27.lut_mask = 64'h00000000F0F00F0F;
defparam fp_functions_0_aadd_2_a27.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_0_a27(
	.dataa(gnd),
	.datab(gnd),
	.datac(!b[26]),
	.datad(!a[26]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_0_a32_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fp_functions_0_aadd_0_a27_cout),
	.shareout());
defparam fp_functions_0_aadd_0_a27.extended_lut = "off";
defparam fp_functions_0_aadd_0_a27.lut_mask = 64'h0000000000F0F00F;
defparam fp_functions_0_aadd_0_a27.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_3_a27(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aadd_1_a6_sumout),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_3_a32_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fp_functions_0_aadd_3_a27_cout),
	.shareout());
defparam fp_functions_0_aadd_3_a27.extended_lut = "off";
defparam fp_functions_0_aadd_3_a27.lut_mask = 64'h0000000000000F0F;
defparam fp_functions_0_aadd_3_a27.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_2_a32(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aadd_1_a1_sumout),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_2_a37_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fp_functions_0_aadd_2_a32_cout),
	.shareout());
defparam fp_functions_0_aadd_2_a32.extended_lut = "off";
defparam fp_functions_0_aadd_2_a32.lut_mask = 64'h00000000F0F00F0F;
defparam fp_functions_0_aadd_2_a32.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_0_a32(
	.dataa(gnd),
	.datab(gnd),
	.datac(!b[25]),
	.datad(!a[25]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_0_a37_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fp_functions_0_aadd_0_a32_cout),
	.shareout());
defparam fp_functions_0_aadd_0_a32.extended_lut = "off";
defparam fp_functions_0_aadd_0_a32.lut_mask = 64'h0000000000F0F00F;
defparam fp_functions_0_aadd_0_a32.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_3_a32(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aadd_1_a1_sumout),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_3_a37_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fp_functions_0_aadd_3_a32_cout),
	.shareout());
defparam fp_functions_0_aadd_3_a32.extended_lut = "off";
defparam fp_functions_0_aadd_3_a32.lut_mask = 64'h000000000F0FF0F0;
defparam fp_functions_0_aadd_3_a32.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_2_a37(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aadd_1_a21_sumout),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_2_a42_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fp_functions_0_aadd_2_a37_cout),
	.shareout());
defparam fp_functions_0_aadd_2_a37.extended_lut = "off";
defparam fp_functions_0_aadd_2_a37.lut_mask = 64'h000000000000F0F0;
defparam fp_functions_0_aadd_2_a37.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_0_a37(
	.dataa(gnd),
	.datab(gnd),
	.datac(!b[24]),
	.datad(!a[24]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_0_a42_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fp_functions_0_aadd_0_a37_cout),
	.shareout());
defparam fp_functions_0_aadd_0_a37.extended_lut = "off";
defparam fp_functions_0_aadd_0_a37.lut_mask = 64'h0000000000F0F00F;
defparam fp_functions_0_aadd_0_a37.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_3_a37(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aadd_1_a21_sumout),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_3_a42_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fp_functions_0_aadd_3_a37_cout),
	.shareout());
defparam fp_functions_0_aadd_3_a37.extended_lut = "off";
defparam fp_functions_0_aadd_3_a37.lut_mask = 64'h000000000F0FF0F0;
defparam fp_functions_0_aadd_3_a37.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_2_a42(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aadd_1_a16_sumout),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_2_a47_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fp_functions_0_aadd_2_a42_cout),
	.shareout());
defparam fp_functions_0_aadd_2_a42.extended_lut = "off";
defparam fp_functions_0_aadd_2_a42.lut_mask = 64'h000000000000F0F0;
defparam fp_functions_0_aadd_2_a42.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_0_a42(
	.dataa(gnd),
	.datab(gnd),
	.datac(!b[23]),
	.datad(!a[23]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_0_a47_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fp_functions_0_aadd_0_a42_cout),
	.shareout());
defparam fp_functions_0_aadd_0_a42.extended_lut = "off";
defparam fp_functions_0_aadd_0_a42.lut_mask = 64'h0000000000F0F00F;
defparam fp_functions_0_aadd_0_a42.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_3_a42(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aadd_1_a16_sumout),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_3_a47_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fp_functions_0_aadd_3_a42_cout),
	.shareout());
defparam fp_functions_0_aadd_3_a42.extended_lut = "off";
defparam fp_functions_0_aadd_3_a42.lut_mask = 64'h000000000F0FF0F0;
defparam fp_functions_0_aadd_3_a42.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_2_a47(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aadd_1_a11_sumout),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_2_a52_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fp_functions_0_aadd_2_a47_cout),
	.shareout());
defparam fp_functions_0_aadd_2_a47.extended_lut = "off";
defparam fp_functions_0_aadd_2_a47.lut_mask = 64'h00000000F0F00F0F;
defparam fp_functions_0_aadd_2_a47.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_0_a47(
	.dataa(gnd),
	.datab(gnd),
	.datac(!b[22]),
	.datad(!a[22]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_0_a52_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fp_functions_0_aadd_0_a47_cout),
	.shareout());
defparam fp_functions_0_aadd_0_a47.extended_lut = "off";
defparam fp_functions_0_aadd_0_a47.lut_mask = 64'h0000000000F0F00F;
defparam fp_functions_0_aadd_0_a47.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_3_a47(
	.dataa(gnd),
	.datab(gnd),
	.datac(!fp_functions_0_aadd_1_a11_sumout),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fp_functions_0_aadd_3_a47_cout),
	.shareout());
defparam fp_functions_0_aadd_3_a47.extended_lut = "off";
defparam fp_functions_0_aadd_3_a47.lut_mask = 64'h000000000F0FF0F0;
defparam fp_functions_0_aadd_3_a47.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_2_a52(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fp_functions_0_aadd_2_a52_cout),
	.shareout());
defparam fp_functions_0_aadd_2_a52.extended_lut = "off";
defparam fp_functions_0_aadd_2_a52.lut_mask = 64'h00000000FFFF0000;
defparam fp_functions_0_aadd_2_a52.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_0_a52(
	.dataa(gnd),
	.datab(gnd),
	.datac(!b[21]),
	.datad(!a[21]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_0_a57_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fp_functions_0_aadd_0_a52_cout),
	.shareout());
defparam fp_functions_0_aadd_0_a52.extended_lut = "off";
defparam fp_functions_0_aadd_0_a52.lut_mask = 64'h0000000000F0F00F;
defparam fp_functions_0_aadd_0_a52.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_0_a57(
	.dataa(gnd),
	.datab(gnd),
	.datac(!b[20]),
	.datad(!a[20]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_0_a62_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fp_functions_0_aadd_0_a57_cout),
	.shareout());
defparam fp_functions_0_aadd_0_a57.extended_lut = "off";
defparam fp_functions_0_aadd_0_a57.lut_mask = 64'h0000000000F0F00F;
defparam fp_functions_0_aadd_0_a57.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_0_a62(
	.dataa(gnd),
	.datab(gnd),
	.datac(!b[19]),
	.datad(!a[19]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_0_a67_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fp_functions_0_aadd_0_a62_cout),
	.shareout());
defparam fp_functions_0_aadd_0_a62.extended_lut = "off";
defparam fp_functions_0_aadd_0_a62.lut_mask = 64'h0000000000F0F00F;
defparam fp_functions_0_aadd_0_a62.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_0_a67(
	.dataa(gnd),
	.datab(gnd),
	.datac(!b[18]),
	.datad(!a[18]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_0_a72_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fp_functions_0_aadd_0_a67_cout),
	.shareout());
defparam fp_functions_0_aadd_0_a67.extended_lut = "off";
defparam fp_functions_0_aadd_0_a67.lut_mask = 64'h0000000000F0F00F;
defparam fp_functions_0_aadd_0_a67.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_0_a72(
	.dataa(gnd),
	.datab(gnd),
	.datac(!b[17]),
	.datad(!a[17]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_0_a77_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fp_functions_0_aadd_0_a72_cout),
	.shareout());
defparam fp_functions_0_aadd_0_a72.extended_lut = "off";
defparam fp_functions_0_aadd_0_a72.lut_mask = 64'h0000000000F0F00F;
defparam fp_functions_0_aadd_0_a72.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_0_a77(
	.dataa(gnd),
	.datab(gnd),
	.datac(!b[16]),
	.datad(!a[16]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_0_a82_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fp_functions_0_aadd_0_a77_cout),
	.shareout());
defparam fp_functions_0_aadd_0_a77.extended_lut = "off";
defparam fp_functions_0_aadd_0_a77.lut_mask = 64'h0000000000F0F00F;
defparam fp_functions_0_aadd_0_a77.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_0_a82(
	.dataa(gnd),
	.datab(gnd),
	.datac(!b[15]),
	.datad(!a[15]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_0_a87_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fp_functions_0_aadd_0_a82_cout),
	.shareout());
defparam fp_functions_0_aadd_0_a82.extended_lut = "off";
defparam fp_functions_0_aadd_0_a82.lut_mask = 64'h0000000000F0F00F;
defparam fp_functions_0_aadd_0_a82.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_0_a87(
	.dataa(gnd),
	.datab(gnd),
	.datac(!b[14]),
	.datad(!a[14]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_0_a92_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fp_functions_0_aadd_0_a87_cout),
	.shareout());
defparam fp_functions_0_aadd_0_a87.extended_lut = "off";
defparam fp_functions_0_aadd_0_a87.lut_mask = 64'h0000000000F0F00F;
defparam fp_functions_0_aadd_0_a87.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_0_a92(
	.dataa(gnd),
	.datab(gnd),
	.datac(!b[13]),
	.datad(!a[13]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_0_a97_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fp_functions_0_aadd_0_a92_cout),
	.shareout());
defparam fp_functions_0_aadd_0_a92.extended_lut = "off";
defparam fp_functions_0_aadd_0_a92.lut_mask = 64'h0000000000F0F00F;
defparam fp_functions_0_aadd_0_a92.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_0_a97(
	.dataa(gnd),
	.datab(gnd),
	.datac(!b[12]),
	.datad(!a[12]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_0_a102_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fp_functions_0_aadd_0_a97_cout),
	.shareout());
defparam fp_functions_0_aadd_0_a97.extended_lut = "off";
defparam fp_functions_0_aadd_0_a97.lut_mask = 64'h0000000000F0F00F;
defparam fp_functions_0_aadd_0_a97.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_0_a102(
	.dataa(gnd),
	.datab(gnd),
	.datac(!b[11]),
	.datad(!a[11]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_0_a107_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fp_functions_0_aadd_0_a102_cout),
	.shareout());
defparam fp_functions_0_aadd_0_a102.extended_lut = "off";
defparam fp_functions_0_aadd_0_a102.lut_mask = 64'h0000000000F0F00F;
defparam fp_functions_0_aadd_0_a102.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_0_a107(
	.dataa(gnd),
	.datab(gnd),
	.datac(!b[10]),
	.datad(!a[10]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_0_a112_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fp_functions_0_aadd_0_a107_cout),
	.shareout());
defparam fp_functions_0_aadd_0_a107.extended_lut = "off";
defparam fp_functions_0_aadd_0_a107.lut_mask = 64'h0000000000F0F00F;
defparam fp_functions_0_aadd_0_a107.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_0_a112(
	.dataa(gnd),
	.datab(gnd),
	.datac(!b[9]),
	.datad(!a[9]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_0_a117_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fp_functions_0_aadd_0_a112_cout),
	.shareout());
defparam fp_functions_0_aadd_0_a112.extended_lut = "off";
defparam fp_functions_0_aadd_0_a112.lut_mask = 64'h0000000000F0F00F;
defparam fp_functions_0_aadd_0_a112.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_0_a117(
	.dataa(gnd),
	.datab(gnd),
	.datac(!b[8]),
	.datad(!a[8]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_0_a122_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fp_functions_0_aadd_0_a117_cout),
	.shareout());
defparam fp_functions_0_aadd_0_a117.extended_lut = "off";
defparam fp_functions_0_aadd_0_a117.lut_mask = 64'h0000000000F0F00F;
defparam fp_functions_0_aadd_0_a117.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_0_a122(
	.dataa(gnd),
	.datab(gnd),
	.datac(!b[7]),
	.datad(!a[7]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_0_a127_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fp_functions_0_aadd_0_a122_cout),
	.shareout());
defparam fp_functions_0_aadd_0_a122.extended_lut = "off";
defparam fp_functions_0_aadd_0_a122.lut_mask = 64'h0000000000F0F00F;
defparam fp_functions_0_aadd_0_a122.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_0_a127(
	.dataa(gnd),
	.datab(gnd),
	.datac(!b[6]),
	.datad(!a[6]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_0_a132_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fp_functions_0_aadd_0_a127_cout),
	.shareout());
defparam fp_functions_0_aadd_0_a127.extended_lut = "off";
defparam fp_functions_0_aadd_0_a127.lut_mask = 64'h0000000000F0F00F;
defparam fp_functions_0_aadd_0_a127.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_0_a132(
	.dataa(gnd),
	.datab(gnd),
	.datac(!b[5]),
	.datad(!a[5]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_0_a137_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fp_functions_0_aadd_0_a132_cout),
	.shareout());
defparam fp_functions_0_aadd_0_a132.extended_lut = "off";
defparam fp_functions_0_aadd_0_a132.lut_mask = 64'h0000000000F0F00F;
defparam fp_functions_0_aadd_0_a132.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_0_a137(
	.dataa(gnd),
	.datab(gnd),
	.datac(!b[4]),
	.datad(!a[4]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_0_a142_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fp_functions_0_aadd_0_a137_cout),
	.shareout());
defparam fp_functions_0_aadd_0_a137.extended_lut = "off";
defparam fp_functions_0_aadd_0_a137.lut_mask = 64'h0000000000F0F00F;
defparam fp_functions_0_aadd_0_a137.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_0_a142(
	.dataa(gnd),
	.datab(gnd),
	.datac(!b[3]),
	.datad(!a[3]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_0_a147_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fp_functions_0_aadd_0_a142_cout),
	.shareout());
defparam fp_functions_0_aadd_0_a142.extended_lut = "off";
defparam fp_functions_0_aadd_0_a142.lut_mask = 64'h0000000000F0F00F;
defparam fp_functions_0_aadd_0_a142.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_0_a147(
	.dataa(gnd),
	.datab(gnd),
	.datac(!b[2]),
	.datad(!a[2]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_0_a152_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fp_functions_0_aadd_0_a147_cout),
	.shareout());
defparam fp_functions_0_aadd_0_a147.extended_lut = "off";
defparam fp_functions_0_aadd_0_a147.lut_mask = 64'h0000000000F0F00F;
defparam fp_functions_0_aadd_0_a147.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_0_a152(
	.dataa(gnd),
	.datab(gnd),
	.datac(!b[1]),
	.datad(!a[1]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_0_a157_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fp_functions_0_aadd_0_a152_cout),
	.shareout());
defparam fp_functions_0_aadd_0_a152.extended_lut = "off";
defparam fp_functions_0_aadd_0_a152.lut_mask = 64'h0000000000F0F00F;
defparam fp_functions_0_aadd_0_a152.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_0_a157(
	.dataa(gnd),
	.datab(gnd),
	.datac(!b[0]),
	.datad(!a[0]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(fp_functions_0_aadd_0_a162_cout),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fp_functions_0_aadd_0_a157_cout),
	.shareout());
defparam fp_functions_0_aadd_0_a157.extended_lut = "off";
defparam fp_functions_0_aadd_0_a157.lut_mask = 64'h0000000000F0F00F;
defparam fp_functions_0_aadd_0_a157.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aadd_0_a162(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(fp_functions_0_aadd_0_a162_cout),
	.shareout());
defparam fp_functions_0_aadd_0_a162.extended_lut = "off";
defparam fp_functions_0_aadd_0_a162.lut_mask = 64'h00000000FFFF0000;
defparam fp_functions_0_aadd_0_a162.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_areduce_nor_7_a3(
	.dataa(!fp_functions_0_areduce_nor_7_a2_combout),
	.datab(!fp_functions_0_areduce_nor_7_a1_combout),
	.datac(!fp_functions_0_areduce_nor_7_a0_combout),
	.datad(!a[25]),
	.datae(!fp_functions_0_aexp_bSig_uid35_fpAddTest_b_a3_a_a0_combout),
	.dataf(!fp_functions_0_areduce_nor_7_a0_combout),
	.datag(!b[25]),
	.datah(!fp_functions_0_aadd_0_a1_sumout),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_areduce_nor_7_a3_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_areduce_nor_7_a3.extended_lut = "on";
defparam fp_functions_0_areduce_nor_7_a3.lut_mask = 64'h0000008000000080;
defparam fp_functions_0_areduce_nor_7_a3.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai1783_a34(
	.dataa(!fp_functions_0_aadd_1_a1_sumout),
	.datab(!fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a2_a_a1_combout),
	.datac(!fp_functions_0_aMux_58_a1_combout),
	.datad(!fp_functions_0_aMux_58_a0_combout),
	.datae(!fp_functions_0_aadd_1_a16_sumout),
	.dataf(!fp_functions_0_aMux_54_a1_combout),
	.datag(!fp_functions_0_aMux_2_a25_combout),
	.datah(!fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a13_a_a2_combout),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai1783_a34_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai1783_a34.extended_lut = "on";
defparam fp_functions_0_ai1783_a34.lut_mask = 64'h0C0C0C3F084C084C;
defparam fp_functions_0_ai1783_a34.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai1783_a39(
	.dataa(!fp_functions_0_aadd_1_a1_sumout),
	.datab(!fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a2_a_a1_combout),
	.datac(!fp_functions_0_aMux_59_a6_combout),
	.datad(!fp_functions_0_aMux_59_a5_combout),
	.datae(!fp_functions_0_aadd_1_a16_sumout),
	.dataf(!fp_functions_0_aMux_55_a1_combout),
	.datag(!fp_functions_0_aMux_2_a10_combout),
	.datah(!fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a13_a_a2_combout),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai1783_a39_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai1783_a39.extended_lut = "on";
defparam fp_functions_0_ai1783_a39.lut_mask = 64'h0C0C0C3F084C084C;
defparam fp_functions_0_ai1783_a39.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_55_a1(
	.dataa(!fp_functions_0_aadd_1_a1_sumout),
	.datab(!fp_functions_0_aMux_2_a13_combout),
	.datac(gnd),
	.datad(!fp_functions_0_aMux_2_a11_combout),
	.datae(!fp_functions_0_aadd_1_a16_sumout),
	.dataf(!fp_functions_0_aMux_2_a3_combout),
	.datag(!fp_functions_0_aMux_2_a2_combout),
	.datah(!fp_functions_0_aadd_1_a21_sumout),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_55_a1_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_55_a1.extended_lut = "on";
defparam fp_functions_0_aMux_55_a1.lut_mask = 64'h00AA0A0A222200AA;
defparam fp_functions_0_aMux_55_a1.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai1783_a44(
	.dataa(!fp_functions_0_aMux_2_a8_combout),
	.datab(!fp_functions_0_aadd_1_a16_sumout),
	.datac(!fp_functions_0_aMux_2_a10_combout),
	.datad(!fp_functions_0_areduce_nor_0_acombout),
	.datae(!fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a13_a_a2_combout),
	.dataf(!fp_functions_0_aMux_53_a1_combout),
	.datag(!fp_functions_0_ai1783_a19_combout),
	.datah(!fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a2_a_a1_combout),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai1783_a44_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai1783_a44.extended_lut = "on";
defparam fp_functions_0_ai1783_a44.lut_mask = 64'h0F0F00FF0C1D0000;
defparam fp_functions_0_ai1783_a44.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai1783_a49(
	.dataa(!fp_functions_0_aMux_23_a0_combout),
	.datab(!fp_functions_0_aadd_1_a16_sumout),
	.datac(!fp_functions_0_areduce_nor_0_acombout),
	.datad(!fp_functions_0_aMux_23_a1_combout),
	.datae(!fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a13_a_a2_combout),
	.dataf(!fp_functions_0_ai1783_a18_combout),
	.datag(!fp_functions_0_aMux_52_a0_combout),
	.datah(!fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a2_a_a1_combout),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai1783_a49_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai1783_a49.extended_lut = "on";
defparam fp_functions_0_ai1783_a49.lut_mask = 64'h00FF0F0F04070000;
defparam fp_functions_0_ai1783_a49.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_204_a0(
	.dataa(!fp_functions_0_aregInputs_uid118_fpAddTest_delay_adelay_signals_a0_a_a0_a_aq),
	.datab(!fp_functions_0_aredist16_excZ_aSig_uid16_uid23_fpAddTest_q_1_q_a0_a_aq),
	.datac(!fp_functions_0_aredist14_excZ_bSig_uid17_uid37_fpAddTest_q_3_q_a0_a_aq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_204_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_204_a0.extended_lut = "off";
defparam fp_functions_0_aMux_204_a0.lut_mask = 64'h4242424242424242;
defparam fp_functions_0_aMux_204_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_236_a0(
	.dataa(!fp_functions_0_aredist4_effSub_uid52_fpAddTest_q_2_q_a0_a_aq),
	.datab(!fp_functions_0_aredist15_excI_aSig_uid27_fpAddTest_q_1_q_a0_a_aq),
	.datac(!fp_functions_0_aredist10_excI_bSig_uid41_fpAddTest_q_1_q_a0_a_aq),
	.datad(!fp_functions_0_aexcN_bSig_uid42_fpAddTest_delay_adelay_signals_a0_a_a0_a_aq),
	.datae(!fp_functions_0_aexcN_aSig_uid28_fpAddTest_delay_adelay_signals_a0_a_a0_a_aq),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_236_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_236_a0.extended_lut = "off";
defparam fp_functions_0_aMux_236_a0.lut_mask = 64'hFE000000FE000000;
defparam fp_functions_0_aMux_236_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_areduce_nor_15_a0(
	.dataa(!fp_functions_0_aadd_7_a11_sumout),
	.datab(!fp_functions_0_aadd_7_a16_sumout),
	.datac(!fp_functions_0_aadd_7_a21_sumout),
	.datad(!fp_functions_0_aadd_7_a26_sumout),
	.datae(!fp_functions_0_aadd_7_a31_sumout),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_areduce_nor_15_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_areduce_nor_15_a0.extended_lut = "off";
defparam fp_functions_0_areduce_nor_15_a0.lut_mask = 64'h8000000080000000;
defparam fp_functions_0_areduce_nor_15_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aexcRZeroVInC_uid119_fpAddTest_q_a3_a(
	.dataa(!fp_functions_0_aadd_7_a6_sumout),
	.datab(!fp_functions_0_areduce_nor_15_a0_combout),
	.datac(!fp_functions_0_aadd_7_a36_sumout),
	.datad(!fp_functions_0_aadd_7_a41_sumout),
	.datae(!fp_functions_0_aadd_7_a46_sumout),
	.dataf(!fp_functions_0_aadd_7_a51_sumout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aexcRZeroVInC_uid119_fpAddTest_q_a3_a_acombout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aexcRZeroVInC_uid119_fpAddTest_q_a3_a.extended_lut = "off";
defparam fp_functions_0_aexcRZeroVInC_uid119_fpAddTest_q_a3_a.lut_mask = 64'hDFFFFFFF00000000;
defparam fp_functions_0_aexcRZeroVInC_uid119_fpAddTest_q_a3_a.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_204_a1(
	.dataa(!fp_functions_0_aredist16_excZ_aSig_uid16_uid23_fpAddTest_q_1_q_a0_a_aq),
	.datab(!fp_functions_0_aredist14_excZ_bSig_uid17_uid37_fpAddTest_q_3_q_a0_a_aq),
	.datac(!fp_functions_0_aregInputs_uid118_fpAddTest_delay_adelay_signals_a0_a_a0_a_aq),
	.datad(!fp_functions_0_aexcRZeroVInC_uid119_fpAddTest_q_a3_a_acombout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_204_a1_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_204_a1.extended_lut = "off";
defparam fp_functions_0_aMux_204_a1.lut_mask = 64'h1810181018101810;
defparam fp_functions_0_aMux_204_a1.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aexcRInfVInC_uid122_fpAddTest_q_a5_a_a0(
	.dataa(!fp_functions_0_aadd_7_a11_sumout),
	.datab(!fp_functions_0_aadd_7_a16_sumout),
	.datac(!fp_functions_0_aadd_7_a21_sumout),
	.datad(!fp_functions_0_aadd_7_a26_sumout),
	.datae(!fp_functions_0_aadd_7_a31_sumout),
	.dataf(!fp_functions_0_aadd_7_a6_sumout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aexcRInfVInC_uid122_fpAddTest_q_a5_a_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aexcRInfVInC_uid122_fpAddTest_q_a5_a_a0.extended_lut = "off";
defparam fp_functions_0_aexcRInfVInC_uid122_fpAddTest_q_a5_a_a0.lut_mask = 64'h0000000000000001;
defparam fp_functions_0_aexcRInfVInC_uid122_fpAddTest_q_a5_a_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aexcRInfVInC_uid122_fpAddTest_q_a5_a_a1(
	.dataa(!fp_functions_0_aregInputs_uid118_fpAddTest_delay_adelay_signals_a0_a_a0_a_aq),
	.datab(!fp_functions_0_aadd_7_a36_sumout),
	.datac(!fp_functions_0_aexcRInfVInC_uid122_fpAddTest_q_a5_a_a0_combout),
	.datad(!fp_functions_0_aadd_7_a41_sumout),
	.datae(!fp_functions_0_aadd_7_a46_sumout),
	.dataf(!fp_functions_0_aadd_7_a51_sumout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aexcRInfVInC_uid122_fpAddTest_q_a5_a_a1_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aexcRInfVInC_uid122_fpAddTest_q_a5_a_a1.extended_lut = "off";
defparam fp_functions_0_aexcRInfVInC_uid122_fpAddTest_q_a5_a_a1.lut_mask = 64'h0001555500000000;
defparam fp_functions_0_aexcRInfVInC_uid122_fpAddTest_q_a5_a_a1.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_203_a2(
	.dataa(!fp_functions_0_aredist4_effSub_uid52_fpAddTest_q_2_q_a0_a_aq),
	.datab(!fp_functions_0_aredist15_excI_aSig_uid27_fpAddTest_q_1_q_a0_a_aq),
	.datac(!fp_functions_0_aredist10_excI_bSig_uid41_fpAddTest_q_1_q_a0_a_aq),
	.datad(!fp_functions_0_aexcRInfVInC_uid122_fpAddTest_q_a5_a_a1_combout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_203_a2_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_203_a2.extended_lut = "off";
defparam fp_functions_0_aMux_203_a2.lut_mask = 64'h3E803E803E803E80;
defparam fp_functions_0_aMux_203_a2.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_237_a2(
	.dataa(!fp_functions_0_aredist2_aMinusA_uid87_fpAddTest_q_1_q_a0_a_aq),
	.datab(!fp_functions_0_aMux_204_a0_combout),
	.datac(!fp_functions_0_aMux_236_a0_combout),
	.datad(!fp_functions_0_aadd_7_a1_sumout),
	.datae(!fp_functions_0_aMux_204_a1_combout),
	.dataf(!fp_functions_0_aMux_203_a2_combout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_237_a2_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_237_a2.extended_lut = "off";
defparam fp_functions_0_aMux_237_a2.lut_mask = 64'hF0FEF0F4F0F0F0F0;
defparam fp_functions_0_aMux_237_a2.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_236_a1(
	.dataa(!fp_functions_0_aredist2_aMinusA_uid87_fpAddTest_q_1_q_a0_a_aq),
	.datab(!fp_functions_0_aMux_204_a0_combout),
	.datac(!fp_functions_0_aMux_236_a0_combout),
	.datad(!fp_functions_0_aadd_7_a56_sumout),
	.datae(!fp_functions_0_aMux_204_a1_combout),
	.dataf(!fp_functions_0_aMux_203_a2_combout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_236_a1_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_236_a1.extended_lut = "off";
defparam fp_functions_0_aMux_236_a1.lut_mask = 64'h000E000400000000;
defparam fp_functions_0_aMux_236_a1.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_235_a0(
	.dataa(!fp_functions_0_aredist2_aMinusA_uid87_fpAddTest_q_1_q_a0_a_aq),
	.datab(!fp_functions_0_aMux_204_a0_combout),
	.datac(!fp_functions_0_aMux_236_a0_combout),
	.datad(!fp_functions_0_aadd_7_a61_sumout),
	.datae(!fp_functions_0_aMux_204_a1_combout),
	.dataf(!fp_functions_0_aMux_203_a2_combout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_235_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_235_a0.extended_lut = "off";
defparam fp_functions_0_aMux_235_a0.lut_mask = 64'h000E000400000000;
defparam fp_functions_0_aMux_235_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_234_a0(
	.dataa(!fp_functions_0_aredist2_aMinusA_uid87_fpAddTest_q_1_q_a0_a_aq),
	.datab(!fp_functions_0_aMux_204_a0_combout),
	.datac(!fp_functions_0_aMux_236_a0_combout),
	.datad(!fp_functions_0_aadd_7_a66_sumout),
	.datae(!fp_functions_0_aMux_204_a1_combout),
	.dataf(!fp_functions_0_aMux_203_a2_combout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_234_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_234_a0.extended_lut = "off";
defparam fp_functions_0_aMux_234_a0.lut_mask = 64'h000E000400000000;
defparam fp_functions_0_aMux_234_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_233_a0(
	.dataa(!fp_functions_0_aredist2_aMinusA_uid87_fpAddTest_q_1_q_a0_a_aq),
	.datab(!fp_functions_0_aMux_204_a0_combout),
	.datac(!fp_functions_0_aMux_236_a0_combout),
	.datad(!fp_functions_0_aadd_7_a71_sumout),
	.datae(!fp_functions_0_aMux_204_a1_combout),
	.dataf(!fp_functions_0_aMux_203_a2_combout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_233_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_233_a0.extended_lut = "off";
defparam fp_functions_0_aMux_233_a0.lut_mask = 64'h000E000400000000;
defparam fp_functions_0_aMux_233_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_232_a0(
	.dataa(!fp_functions_0_aredist2_aMinusA_uid87_fpAddTest_q_1_q_a0_a_aq),
	.datab(!fp_functions_0_aMux_204_a0_combout),
	.datac(!fp_functions_0_aMux_236_a0_combout),
	.datad(!fp_functions_0_aadd_7_a76_sumout),
	.datae(!fp_functions_0_aMux_204_a1_combout),
	.dataf(!fp_functions_0_aMux_203_a2_combout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_232_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_232_a0.extended_lut = "off";
defparam fp_functions_0_aMux_232_a0.lut_mask = 64'h000E000400000000;
defparam fp_functions_0_aMux_232_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_231_a0(
	.dataa(!fp_functions_0_aredist2_aMinusA_uid87_fpAddTest_q_1_q_a0_a_aq),
	.datab(!fp_functions_0_aMux_204_a0_combout),
	.datac(!fp_functions_0_aMux_236_a0_combout),
	.datad(!fp_functions_0_aadd_7_a81_sumout),
	.datae(!fp_functions_0_aMux_204_a1_combout),
	.dataf(!fp_functions_0_aMux_203_a2_combout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_231_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_231_a0.extended_lut = "off";
defparam fp_functions_0_aMux_231_a0.lut_mask = 64'h000E000400000000;
defparam fp_functions_0_aMux_231_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_230_a0(
	.dataa(!fp_functions_0_aredist2_aMinusA_uid87_fpAddTest_q_1_q_a0_a_aq),
	.datab(!fp_functions_0_aMux_204_a0_combout),
	.datac(!fp_functions_0_aMux_236_a0_combout),
	.datad(!fp_functions_0_aadd_7_a86_sumout),
	.datae(!fp_functions_0_aMux_204_a1_combout),
	.dataf(!fp_functions_0_aMux_203_a2_combout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_230_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_230_a0.extended_lut = "off";
defparam fp_functions_0_aMux_230_a0.lut_mask = 64'h000E000400000000;
defparam fp_functions_0_aMux_230_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_229_a0(
	.dataa(!fp_functions_0_aredist2_aMinusA_uid87_fpAddTest_q_1_q_a0_a_aq),
	.datab(!fp_functions_0_aMux_204_a0_combout),
	.datac(!fp_functions_0_aMux_236_a0_combout),
	.datad(!fp_functions_0_aadd_7_a91_sumout),
	.datae(!fp_functions_0_aMux_204_a1_combout),
	.dataf(!fp_functions_0_aMux_203_a2_combout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_229_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_229_a0.extended_lut = "off";
defparam fp_functions_0_aMux_229_a0.lut_mask = 64'h000E000400000000;
defparam fp_functions_0_aMux_229_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_228_a0(
	.dataa(!fp_functions_0_aredist2_aMinusA_uid87_fpAddTest_q_1_q_a0_a_aq),
	.datab(!fp_functions_0_aMux_204_a0_combout),
	.datac(!fp_functions_0_aMux_236_a0_combout),
	.datad(!fp_functions_0_aadd_7_a96_sumout),
	.datae(!fp_functions_0_aMux_204_a1_combout),
	.dataf(!fp_functions_0_aMux_203_a2_combout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_228_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_228_a0.extended_lut = "off";
defparam fp_functions_0_aMux_228_a0.lut_mask = 64'h000E000400000000;
defparam fp_functions_0_aMux_228_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_227_a0(
	.dataa(!fp_functions_0_aredist2_aMinusA_uid87_fpAddTest_q_1_q_a0_a_aq),
	.datab(!fp_functions_0_aMux_204_a0_combout),
	.datac(!fp_functions_0_aMux_236_a0_combout),
	.datad(!fp_functions_0_aadd_7_a101_sumout),
	.datae(!fp_functions_0_aMux_204_a1_combout),
	.dataf(!fp_functions_0_aMux_203_a2_combout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_227_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_227_a0.extended_lut = "off";
defparam fp_functions_0_aMux_227_a0.lut_mask = 64'h000E000400000000;
defparam fp_functions_0_aMux_227_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_226_a0(
	.dataa(!fp_functions_0_aredist2_aMinusA_uid87_fpAddTest_q_1_q_a0_a_aq),
	.datab(!fp_functions_0_aMux_204_a0_combout),
	.datac(!fp_functions_0_aMux_236_a0_combout),
	.datad(!fp_functions_0_aadd_7_a106_sumout),
	.datae(!fp_functions_0_aMux_204_a1_combout),
	.dataf(!fp_functions_0_aMux_203_a2_combout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_226_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_226_a0.extended_lut = "off";
defparam fp_functions_0_aMux_226_a0.lut_mask = 64'h000E000400000000;
defparam fp_functions_0_aMux_226_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_225_a0(
	.dataa(!fp_functions_0_aredist2_aMinusA_uid87_fpAddTest_q_1_q_a0_a_aq),
	.datab(!fp_functions_0_aMux_204_a0_combout),
	.datac(!fp_functions_0_aMux_236_a0_combout),
	.datad(!fp_functions_0_aadd_7_a111_sumout),
	.datae(!fp_functions_0_aMux_204_a1_combout),
	.dataf(!fp_functions_0_aMux_203_a2_combout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_225_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_225_a0.extended_lut = "off";
defparam fp_functions_0_aMux_225_a0.lut_mask = 64'h000E000400000000;
defparam fp_functions_0_aMux_225_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_224_a0(
	.dataa(!fp_functions_0_aredist2_aMinusA_uid87_fpAddTest_q_1_q_a0_a_aq),
	.datab(!fp_functions_0_aMux_204_a0_combout),
	.datac(!fp_functions_0_aMux_236_a0_combout),
	.datad(!fp_functions_0_aadd_7_a116_sumout),
	.datae(!fp_functions_0_aMux_204_a1_combout),
	.dataf(!fp_functions_0_aMux_203_a2_combout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_224_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_224_a0.extended_lut = "off";
defparam fp_functions_0_aMux_224_a0.lut_mask = 64'h000E000400000000;
defparam fp_functions_0_aMux_224_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_223_a0(
	.dataa(!fp_functions_0_aredist2_aMinusA_uid87_fpAddTest_q_1_q_a0_a_aq),
	.datab(!fp_functions_0_aMux_204_a0_combout),
	.datac(!fp_functions_0_aMux_236_a0_combout),
	.datad(!fp_functions_0_aadd_7_a121_sumout),
	.datae(!fp_functions_0_aMux_204_a1_combout),
	.dataf(!fp_functions_0_aMux_203_a2_combout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_223_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_223_a0.extended_lut = "off";
defparam fp_functions_0_aMux_223_a0.lut_mask = 64'h000E000400000000;
defparam fp_functions_0_aMux_223_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_222_a0(
	.dataa(!fp_functions_0_aredist2_aMinusA_uid87_fpAddTest_q_1_q_a0_a_aq),
	.datab(!fp_functions_0_aMux_204_a0_combout),
	.datac(!fp_functions_0_aMux_236_a0_combout),
	.datad(!fp_functions_0_aadd_7_a126_sumout),
	.datae(!fp_functions_0_aMux_204_a1_combout),
	.dataf(!fp_functions_0_aMux_203_a2_combout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_222_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_222_a0.extended_lut = "off";
defparam fp_functions_0_aMux_222_a0.lut_mask = 64'h000E000400000000;
defparam fp_functions_0_aMux_222_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_221_a0(
	.dataa(!fp_functions_0_aredist2_aMinusA_uid87_fpAddTest_q_1_q_a0_a_aq),
	.datab(!fp_functions_0_aMux_204_a0_combout),
	.datac(!fp_functions_0_aMux_236_a0_combout),
	.datad(!fp_functions_0_aadd_7_a131_sumout),
	.datae(!fp_functions_0_aMux_204_a1_combout),
	.dataf(!fp_functions_0_aMux_203_a2_combout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_221_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_221_a0.extended_lut = "off";
defparam fp_functions_0_aMux_221_a0.lut_mask = 64'h000E000400000000;
defparam fp_functions_0_aMux_221_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_220_a0(
	.dataa(!fp_functions_0_aredist2_aMinusA_uid87_fpAddTest_q_1_q_a0_a_aq),
	.datab(!fp_functions_0_aMux_204_a0_combout),
	.datac(!fp_functions_0_aMux_236_a0_combout),
	.datad(!fp_functions_0_aadd_7_a136_sumout),
	.datae(!fp_functions_0_aMux_204_a1_combout),
	.dataf(!fp_functions_0_aMux_203_a2_combout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_220_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_220_a0.extended_lut = "off";
defparam fp_functions_0_aMux_220_a0.lut_mask = 64'h000E000400000000;
defparam fp_functions_0_aMux_220_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_219_a0(
	.dataa(!fp_functions_0_aredist2_aMinusA_uid87_fpAddTest_q_1_q_a0_a_aq),
	.datab(!fp_functions_0_aMux_204_a0_combout),
	.datac(!fp_functions_0_aMux_236_a0_combout),
	.datad(!fp_functions_0_aadd_7_a141_sumout),
	.datae(!fp_functions_0_aMux_204_a1_combout),
	.dataf(!fp_functions_0_aMux_203_a2_combout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_219_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_219_a0.extended_lut = "off";
defparam fp_functions_0_aMux_219_a0.lut_mask = 64'h000E000400000000;
defparam fp_functions_0_aMux_219_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_218_a0(
	.dataa(!fp_functions_0_aredist2_aMinusA_uid87_fpAddTest_q_1_q_a0_a_aq),
	.datab(!fp_functions_0_aMux_204_a0_combout),
	.datac(!fp_functions_0_aMux_236_a0_combout),
	.datad(!fp_functions_0_aadd_7_a146_sumout),
	.datae(!fp_functions_0_aMux_204_a1_combout),
	.dataf(!fp_functions_0_aMux_203_a2_combout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_218_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_218_a0.extended_lut = "off";
defparam fp_functions_0_aMux_218_a0.lut_mask = 64'h000E000400000000;
defparam fp_functions_0_aMux_218_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_217_a0(
	.dataa(!fp_functions_0_aredist2_aMinusA_uid87_fpAddTest_q_1_q_a0_a_aq),
	.datab(!fp_functions_0_aMux_204_a0_combout),
	.datac(!fp_functions_0_aMux_236_a0_combout),
	.datad(!fp_functions_0_aadd_7_a151_sumout),
	.datae(!fp_functions_0_aMux_204_a1_combout),
	.dataf(!fp_functions_0_aMux_203_a2_combout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_217_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_217_a0.extended_lut = "off";
defparam fp_functions_0_aMux_217_a0.lut_mask = 64'h000E000400000000;
defparam fp_functions_0_aMux_217_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_216_a0(
	.dataa(!fp_functions_0_aredist2_aMinusA_uid87_fpAddTest_q_1_q_a0_a_aq),
	.datab(!fp_functions_0_aMux_204_a0_combout),
	.datac(!fp_functions_0_aMux_236_a0_combout),
	.datad(!fp_functions_0_aadd_7_a156_sumout),
	.datae(!fp_functions_0_aMux_204_a1_combout),
	.dataf(!fp_functions_0_aMux_203_a2_combout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_216_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_216_a0.extended_lut = "off";
defparam fp_functions_0_aMux_216_a0.lut_mask = 64'h000E000400000000;
defparam fp_functions_0_aMux_216_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_215_a0(
	.dataa(!fp_functions_0_aredist2_aMinusA_uid87_fpAddTest_q_1_q_a0_a_aq),
	.datab(!fp_functions_0_aMux_204_a0_combout),
	.datac(!fp_functions_0_aMux_236_a0_combout),
	.datad(!fp_functions_0_aadd_7_a161_sumout),
	.datae(!fp_functions_0_aMux_204_a1_combout),
	.dataf(!fp_functions_0_aMux_203_a2_combout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_215_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_215_a0.extended_lut = "off";
defparam fp_functions_0_aMux_215_a0.lut_mask = 64'h000E000400000000;
defparam fp_functions_0_aMux_215_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_214_a2(
	.dataa(!fp_functions_0_aredist2_aMinusA_uid87_fpAddTest_q_1_q_a0_a_aq),
	.datab(!fp_functions_0_aMux_204_a0_combout),
	.datac(!fp_functions_0_aMux_236_a0_combout),
	.datad(!fp_functions_0_aadd_7_a11_sumout),
	.datae(!fp_functions_0_aMux_204_a1_combout),
	.dataf(!fp_functions_0_aMux_203_a2_combout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_214_a2_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_214_a2.extended_lut = "off";
defparam fp_functions_0_aMux_214_a2.lut_mask = 64'hF0FEF0F4FFFFFFFF;
defparam fp_functions_0_aMux_214_a2.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_213_a2(
	.dataa(!fp_functions_0_aredist2_aMinusA_uid87_fpAddTest_q_1_q_a0_a_aq),
	.datab(!fp_functions_0_aMux_204_a0_combout),
	.datac(!fp_functions_0_aMux_236_a0_combout),
	.datad(!fp_functions_0_aadd_7_a16_sumout),
	.datae(!fp_functions_0_aMux_204_a1_combout),
	.dataf(!fp_functions_0_aMux_203_a2_combout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_213_a2_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_213_a2.extended_lut = "off";
defparam fp_functions_0_aMux_213_a2.lut_mask = 64'hF0FEF0F4FFFFFFFF;
defparam fp_functions_0_aMux_213_a2.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_212_a2(
	.dataa(!fp_functions_0_aredist2_aMinusA_uid87_fpAddTest_q_1_q_a0_a_aq),
	.datab(!fp_functions_0_aMux_204_a0_combout),
	.datac(!fp_functions_0_aMux_236_a0_combout),
	.datad(!fp_functions_0_aadd_7_a21_sumout),
	.datae(!fp_functions_0_aMux_204_a1_combout),
	.dataf(!fp_functions_0_aMux_203_a2_combout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_212_a2_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_212_a2.extended_lut = "off";
defparam fp_functions_0_aMux_212_a2.lut_mask = 64'hF0FEF0F4FFFFFFFF;
defparam fp_functions_0_aMux_212_a2.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_211_a2(
	.dataa(!fp_functions_0_aredist2_aMinusA_uid87_fpAddTest_q_1_q_a0_a_aq),
	.datab(!fp_functions_0_aMux_204_a0_combout),
	.datac(!fp_functions_0_aMux_236_a0_combout),
	.datad(!fp_functions_0_aadd_7_a26_sumout),
	.datae(!fp_functions_0_aMux_204_a1_combout),
	.dataf(!fp_functions_0_aMux_203_a2_combout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_211_a2_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_211_a2.extended_lut = "off";
defparam fp_functions_0_aMux_211_a2.lut_mask = 64'hF0FEF0F4FFFFFFFF;
defparam fp_functions_0_aMux_211_a2.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_210_a2(
	.dataa(!fp_functions_0_aredist2_aMinusA_uid87_fpAddTest_q_1_q_a0_a_aq),
	.datab(!fp_functions_0_aMux_204_a0_combout),
	.datac(!fp_functions_0_aMux_236_a0_combout),
	.datad(!fp_functions_0_aadd_7_a31_sumout),
	.datae(!fp_functions_0_aMux_204_a1_combout),
	.dataf(!fp_functions_0_aMux_203_a2_combout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_210_a2_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_210_a2.extended_lut = "off";
defparam fp_functions_0_aMux_210_a2.lut_mask = 64'hF0FEF0F4FFFFFFFF;
defparam fp_functions_0_aMux_210_a2.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_209_a2(
	.dataa(!fp_functions_0_aredist2_aMinusA_uid87_fpAddTest_q_1_q_a0_a_aq),
	.datab(!fp_functions_0_aMux_204_a0_combout),
	.datac(!fp_functions_0_aMux_236_a0_combout),
	.datad(!fp_functions_0_aadd_7_a6_sumout),
	.datae(!fp_functions_0_aMux_204_a1_combout),
	.dataf(!fp_functions_0_aMux_203_a2_combout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_209_a2_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_209_a2.extended_lut = "off";
defparam fp_functions_0_aMux_209_a2.lut_mask = 64'hF0FEF0F4FFFFFFFF;
defparam fp_functions_0_aMux_209_a2.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_208_a2(
	.dataa(!fp_functions_0_aredist2_aMinusA_uid87_fpAddTest_q_1_q_a0_a_aq),
	.datab(!fp_functions_0_aMux_204_a0_combout),
	.datac(!fp_functions_0_aMux_236_a0_combout),
	.datad(!fp_functions_0_aadd_7_a36_sumout),
	.datae(!fp_functions_0_aMux_204_a1_combout),
	.dataf(!fp_functions_0_aMux_203_a2_combout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_208_a2_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_208_a2.extended_lut = "off";
defparam fp_functions_0_aMux_208_a2.lut_mask = 64'hF0FEF0F4FFFFFFFF;
defparam fp_functions_0_aMux_208_a2.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_207_a2(
	.dataa(!fp_functions_0_aredist2_aMinusA_uid87_fpAddTest_q_1_q_a0_a_aq),
	.datab(!fp_functions_0_aMux_204_a0_combout),
	.datac(!fp_functions_0_aMux_236_a0_combout),
	.datad(!fp_functions_0_aadd_7_a41_sumout),
	.datae(!fp_functions_0_aMux_204_a1_combout),
	.dataf(!fp_functions_0_aMux_203_a2_combout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_207_a2_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_207_a2.extended_lut = "off";
defparam fp_functions_0_aMux_207_a2.lut_mask = 64'hF0FEF0F4FFFFFFFF;
defparam fp_functions_0_aMux_207_a2.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aR_uid148_fpAddTest_q_a31_a_a0(
	.dataa(!fp_functions_0_asignRInfRZRReg_uid137_fpAddTest_delay_adelay_signals_a0_a_a0_a_aq),
	.datab(!fp_functions_0_aMux_236_a0_combout),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aR_uid148_fpAddTest_q_a31_a_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aR_uid148_fpAddTest_q_a31_a_a0.extended_lut = "off";
defparam fp_functions_0_aR_uid148_fpAddTest_q_a31_a_a0.lut_mask = 64'h1111111111111111;
defparam fp_functions_0_aR_uid148_fpAddTest_q_a31_a_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_arVStage_uid165_lzCountVal_uid85_fpAddTest_merged_bit_select_b_a2_a_a4(
	.dataa(!fp_functions_0_avStagei_uid157_lzCountVal_uid85_fpAddTest_q_a11_a_aq),
	.datab(!fp_functions_0_avStagei_uid157_lzCountVal_uid85_fpAddTest_q_a10_a_aq),
	.datac(!fp_functions_0_avStagei_uid157_lzCountVal_uid85_fpAddTest_q_a8_a_aq),
	.datad(!fp_functions_0_avStagei_uid157_lzCountVal_uid85_fpAddTest_q_a9_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_arVStage_uid165_lzCountVal_uid85_fpAddTest_merged_bit_select_b_a2_a_a4_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_arVStage_uid165_lzCountVal_uid85_fpAddTest_merged_bit_select_b_a2_a_a4.extended_lut = "off";
defparam fp_functions_0_arVStage_uid165_lzCountVal_uid85_fpAddTest_merged_bit_select_b_a2_a_a4.lut_mask = 64'h8000800080008000;
defparam fp_functions_0_arVStage_uid165_lzCountVal_uid85_fpAddTest_merged_bit_select_b_a2_a_a4.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_arVStage_uid165_lzCountVal_uid85_fpAddTest_merged_bit_select_b_a2_a_a5(
	.dataa(!fp_functions_0_avStagei_uid157_lzCountVal_uid85_fpAddTest_q_a12_a_aq),
	.datab(!fp_functions_0_avStagei_uid157_lzCountVal_uid85_fpAddTest_q_a13_a_aq),
	.datac(!fp_functions_0_arVStage_uid165_lzCountVal_uid85_fpAddTest_merged_bit_select_b_a2_a_a4_combout),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_arVStage_uid165_lzCountVal_uid85_fpAddTest_merged_bit_select_b_a2_a_a5_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_arVStage_uid165_lzCountVal_uid85_fpAddTest_merged_bit_select_b_a2_a_a5.extended_lut = "off";
defparam fp_functions_0_arVStage_uid165_lzCountVal_uid85_fpAddTest_merged_bit_select_b_a2_a_a5.lut_mask = 64'h0808080808080808;
defparam fp_functions_0_arVStage_uid165_lzCountVal_uid85_fpAddTest_merged_bit_select_b_a2_a_a5.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_arVStage_uid165_lzCountVal_uid85_fpAddTest_merged_bit_select_b_a3_a_a6(
	.dataa(!fp_functions_0_avStagei_uid157_lzCountVal_uid85_fpAddTest_q_a15_a_aq),
	.datab(!fp_functions_0_avStagei_uid157_lzCountVal_uid85_fpAddTest_q_a14_a_aq),
	.datac(!fp_functions_0_avStagei_uid157_lzCountVal_uid85_fpAddTest_q_a7_a_aq),
	.datad(!fp_functions_0_arVStage_uid165_lzCountVal_uid85_fpAddTest_merged_bit_select_b_a2_a_a5_combout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_arVStage_uid165_lzCountVal_uid85_fpAddTest_merged_bit_select_b_a3_a_a6_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_arVStage_uid165_lzCountVal_uid85_fpAddTest_merged_bit_select_b_a3_a_a6.extended_lut = "off";
defparam fp_functions_0_arVStage_uid165_lzCountVal_uid85_fpAddTest_merged_bit_select_b_a3_a_a6.lut_mask = 64'hAAA2AAA2AAA2AAA2;
defparam fp_functions_0_arVStage_uid165_lzCountVal_uid85_fpAddTest_merged_bit_select_b_a3_a_a6.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_areduce_nor_6_a0(
	.dataa(!fp_functions_0_avStagei_uid157_lzCountVal_uid85_fpAddTest_q_a15_a_aq),
	.datab(!fp_functions_0_avStagei_uid157_lzCountVal_uid85_fpAddTest_q_a6_a_aq),
	.datac(!fp_functions_0_avStagei_uid157_lzCountVal_uid85_fpAddTest_q_a14_a_aq),
	.datad(!fp_functions_0_arVStage_uid165_lzCountVal_uid85_fpAddTest_merged_bit_select_b_a2_a_a5_combout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_areduce_nor_6_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_areduce_nor_6_a0.extended_lut = "off";
defparam fp_functions_0_areduce_nor_6_a0.lut_mask = 64'hF0D0F0D0F0D0F0D0;
defparam fp_functions_0_areduce_nor_6_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_arVStage_uid165_lzCountVal_uid85_fpAddTest_merged_bit_select_b_a1_a_a7(
	.dataa(!fp_functions_0_avStagei_uid157_lzCountVal_uid85_fpAddTest_q_a15_a_aq),
	.datab(!fp_functions_0_avStagei_uid157_lzCountVal_uid85_fpAddTest_q_a14_a_aq),
	.datac(!fp_functions_0_arVStage_uid165_lzCountVal_uid85_fpAddTest_merged_bit_select_b_a2_a_a4_combout),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_arVStage_uid165_lzCountVal_uid85_fpAddTest_merged_bit_select_b_a1_a_a7_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_arVStage_uid165_lzCountVal_uid85_fpAddTest_merged_bit_select_b_a1_a_a7.extended_lut = "off";
defparam fp_functions_0_arVStage_uid165_lzCountVal_uid85_fpAddTest_merged_bit_select_b_a1_a_a7.lut_mask = 64'h0808080808080808;
defparam fp_functions_0_arVStage_uid165_lzCountVal_uid85_fpAddTest_merged_bit_select_b_a1_a_a7.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_areduce_nor_6_a1(
	.dataa(!fp_functions_0_avStagei_uid157_lzCountVal_uid85_fpAddTest_q_a12_a_aq),
	.datab(!fp_functions_0_avStagei_uid157_lzCountVal_uid85_fpAddTest_q_a13_a_aq),
	.datac(!fp_functions_0_avStagei_uid157_lzCountVal_uid85_fpAddTest_q_a5_a_aq),
	.datad(!fp_functions_0_avStagei_uid157_lzCountVal_uid85_fpAddTest_q_a4_a_aq),
	.datae(!fp_functions_0_arVStage_uid165_lzCountVal_uid85_fpAddTest_merged_bit_select_b_a1_a_a7_combout),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_areduce_nor_6_a1_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_areduce_nor_6_a1.extended_lut = "off";
defparam fp_functions_0_areduce_nor_6_a1.lut_mask = 64'h8888800088888000;
defparam fp_functions_0_areduce_nor_6_a1.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_arVStage_uid171_lzCountVal_uid85_fpAddTest_merged_bit_select_b_a1_a_a2(
	.dataa(!fp_functions_0_avStagei_uid157_lzCountVal_uid85_fpAddTest_q_a3_a_aq),
	.datab(!fp_functions_0_avStagei_uid157_lzCountVal_uid85_fpAddTest_q_a10_a_aq),
	.datac(!fp_functions_0_avStagei_uid157_lzCountVal_uid85_fpAddTest_q_a8_a_aq),
	.datad(!fp_functions_0_avStagei_uid157_lzCountVal_uid85_fpAddTest_q_a9_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_arVStage_uid171_lzCountVal_uid85_fpAddTest_merged_bit_select_b_a1_a_a2_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_arVStage_uid171_lzCountVal_uid85_fpAddTest_merged_bit_select_b_a1_a_a2.extended_lut = "off";
defparam fp_functions_0_arVStage_uid171_lzCountVal_uid85_fpAddTest_merged_bit_select_b_a1_a_a2.lut_mask = 64'h4000400040004000;
defparam fp_functions_0_arVStage_uid171_lzCountVal_uid85_fpAddTest_merged_bit_select_b_a1_a_a2.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_arVStage_uid171_lzCountVal_uid85_fpAddTest_merged_bit_select_b_a1_a_a3(
	.dataa(!fp_functions_0_avStagei_uid157_lzCountVal_uid85_fpAddTest_q_a11_a_aq),
	.datab(!fp_functions_0_arVStage_uid171_lzCountVal_uid85_fpAddTest_merged_bit_select_b_a1_a_a2_combout),
	.datac(!fp_functions_0_areduce_nor_6_a0_combout),
	.datad(!fp_functions_0_areduce_nor_6_a1_combout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_arVStage_uid171_lzCountVal_uid85_fpAddTest_merged_bit_select_b_a1_a_a3_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_arVStage_uid171_lzCountVal_uid85_fpAddTest_merged_bit_select_b_a1_a_a3.extended_lut = "off";
defparam fp_functions_0_arVStage_uid171_lzCountVal_uid85_fpAddTest_merged_bit_select_b_a1_a_a3.lut_mask = 64'h0007000700070007;
defparam fp_functions_0_arVStage_uid171_lzCountVal_uid85_fpAddTest_merged_bit_select_b_a1_a_a3.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_arVStage_uid171_lzCountVal_uid85_fpAddTest_merged_bit_select_b_a0_a_a4(
	.dataa(!fp_functions_0_avStagei_uid157_lzCountVal_uid85_fpAddTest_q_a11_a_aq),
	.datab(!fp_functions_0_avStagei_uid157_lzCountVal_uid85_fpAddTest_q_a8_a_aq),
	.datac(!fp_functions_0_avStagei_uid157_lzCountVal_uid85_fpAddTest_q_a9_a_aq),
	.datad(!fp_functions_0_avStagei_uid157_lzCountVal_uid85_fpAddTest_q_a14_a_aq),
	.datae(!fp_functions_0_avStagei_uid157_lzCountVal_uid85_fpAddTest_q_a2_a_aq),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_arVStage_uid171_lzCountVal_uid85_fpAddTest_merged_bit_select_b_a0_a_a4_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_arVStage_uid171_lzCountVal_uid85_fpAddTest_merged_bit_select_b_a0_a_a4.extended_lut = "off";
defparam fp_functions_0_arVStage_uid171_lzCountVal_uid85_fpAddTest_merged_bit_select_b_a0_a_a4.lut_mask = 64'h0000800000008000;
defparam fp_functions_0_arVStage_uid171_lzCountVal_uid85_fpAddTest_merged_bit_select_b_a0_a_a4.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_arVStage_uid171_lzCountVal_uid85_fpAddTest_merged_bit_select_b_a0_a_a5(
	.dataa(!fp_functions_0_avStagei_uid157_lzCountVal_uid85_fpAddTest_q_a10_a_aq),
	.datab(!fp_functions_0_arVStage_uid171_lzCountVal_uid85_fpAddTest_merged_bit_select_b_a0_a_a4_combout),
	.datac(!fp_functions_0_arVStage_uid165_lzCountVal_uid85_fpAddTest_merged_bit_select_b_a3_a_a6_combout),
	.datad(!fp_functions_0_areduce_nor_6_a1_combout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_arVStage_uid171_lzCountVal_uid85_fpAddTest_merged_bit_select_b_a0_a_a5_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_arVStage_uid171_lzCountVal_uid85_fpAddTest_merged_bit_select_b_a0_a_a5.extended_lut = "off";
defparam fp_functions_0_arVStage_uid171_lzCountVal_uid85_fpAddTest_merged_bit_select_b_a0_a_a5.lut_mask = 64'h0007000700070007;
defparam fp_functions_0_arVStage_uid171_lzCountVal_uid85_fpAddTest_merged_bit_select_b_a0_a_a5.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_areduce_nor_5_a0(
	.dataa(!fp_functions_0_areduce_nor_6_a0_combout),
	.datab(!fp_functions_0_arVStage_uid165_lzCountVal_uid85_fpAddTest_merged_bit_select_b_a3_a_a6_combout),
	.datac(!fp_functions_0_arVStage_uid171_lzCountVal_uid85_fpAddTest_merged_bit_select_b_a1_a_a3_combout),
	.datad(!fp_functions_0_arVStage_uid171_lzCountVal_uid85_fpAddTest_merged_bit_select_b_a0_a_a5_combout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_areduce_nor_5_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_areduce_nor_5_a0.extended_lut = "off";
defparam fp_functions_0_areduce_nor_5_a0.lut_mask = 64'hEFFFEFFFEFFFEFFF;
defparam fp_functions_0_areduce_nor_5_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_arVStage_uid171_lzCountVal_uid85_fpAddTest_merged_bit_select_c_a1_a_a1(
	.dataa(!fp_functions_0_avStagei_uid157_lzCountVal_uid85_fpAddTest_q_a11_a_aq),
	.datab(!fp_functions_0_avStagei_uid157_lzCountVal_uid85_fpAddTest_q_a10_a_aq),
	.datac(!fp_functions_0_avStagei_uid157_lzCountVal_uid85_fpAddTest_q_a8_a_aq),
	.datad(!fp_functions_0_avStagei_uid157_lzCountVal_uid85_fpAddTest_q_a9_a_aq),
	.datae(!fp_functions_0_avStagei_uid157_lzCountVal_uid85_fpAddTest_q_a1_a_aq),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_arVStage_uid171_lzCountVal_uid85_fpAddTest_merged_bit_select_c_a1_a_a1_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_arVStage_uid171_lzCountVal_uid85_fpAddTest_merged_bit_select_c_a1_a_a1.extended_lut = "off";
defparam fp_functions_0_arVStage_uid171_lzCountVal_uid85_fpAddTest_merged_bit_select_c_a1_a_a1.lut_mask = 64'hFF007F00FF007F00;
defparam fp_functions_0_arVStage_uid171_lzCountVal_uid85_fpAddTest_merged_bit_select_c_a1_a_a1.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_arVStage_uid171_lzCountVal_uid85_fpAddTest_merged_bit_select_c_a1_a_a2(
	.dataa(!fp_functions_0_avStagei_uid157_lzCountVal_uid85_fpAddTest_q_a12_a_aq),
	.datab(!fp_functions_0_avStagei_uid157_lzCountVal_uid85_fpAddTest_q_a13_a_aq),
	.datac(!fp_functions_0_avStagei_uid157_lzCountVal_uid85_fpAddTest_q_a5_a_aq),
	.datad(!fp_functions_0_avStagei_uid157_lzCountVal_uid85_fpAddTest_q_a4_a_aq),
	.datae(!fp_functions_0_arVStage_uid165_lzCountVal_uid85_fpAddTest_merged_bit_select_b_a1_a_a7_combout),
	.dataf(!fp_functions_0_arVStage_uid171_lzCountVal_uid85_fpAddTest_merged_bit_select_c_a1_a_a1_combout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_arVStage_uid171_lzCountVal_uid85_fpAddTest_merged_bit_select_c_a1_a_a2_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_arVStage_uid171_lzCountVal_uid85_fpAddTest_merged_bit_select_c_a1_a_a2.extended_lut = "off";
defparam fp_functions_0_arVStage_uid171_lzCountVal_uid85_fpAddTest_merged_bit_select_c_a1_a_a2.lut_mask = 64'h444444C4CCCCC4C4;
defparam fp_functions_0_arVStage_uid171_lzCountVal_uid85_fpAddTest_merged_bit_select_c_a1_a_a2.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_arVStage_uid177_lzCountVal_uid85_fpAddTest_b_a0_a_a0(
	.dataa(!fp_functions_0_areduce_nor_6_a0_combout),
	.datab(!fp_functions_0_arVStage_uid171_lzCountVal_uid85_fpAddTest_merged_bit_select_c_a1_a_a2_combout),
	.datac(!fp_functions_0_arVStage_uid171_lzCountVal_uid85_fpAddTest_merged_bit_select_b_a0_a_a5_combout),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_arVStage_uid177_lzCountVal_uid85_fpAddTest_b_a0_a_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_arVStage_uid177_lzCountVal_uid85_fpAddTest_b_a0_a_a0.extended_lut = "off";
defparam fp_functions_0_arVStage_uid177_lzCountVal_uid85_fpAddTest_b_a0_a_a0.lut_mask = 64'h4040404040404040;
defparam fp_functions_0_arVStage_uid177_lzCountVal_uid85_fpAddTest_b_a0_a_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_arVStage_uid177_lzCountVal_uid85_fpAddTest_b_a0_a_a1(
	.dataa(!fp_functions_0_arVStage_uid165_lzCountVal_uid85_fpAddTest_merged_bit_select_b_a3_a_a6_combout),
	.datab(!fp_functions_0_arVStage_uid171_lzCountVal_uid85_fpAddTest_merged_bit_select_b_a1_a_a3_combout),
	.datac(!fp_functions_0_arVStage_uid177_lzCountVal_uid85_fpAddTest_b_a0_a_a0_combout),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_arVStage_uid177_lzCountVal_uid85_fpAddTest_b_a0_a_a1_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_arVStage_uid177_lzCountVal_uid85_fpAddTest_b_a0_a_a1.extended_lut = "off";
defparam fp_functions_0_arVStage_uid177_lzCountVal_uid85_fpAddTest_b_a0_a_a1.lut_mask = 64'h4040404040404040;
defparam fp_functions_0_arVStage_uid177_lzCountVal_uid85_fpAddTest_b_a0_a_a1.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_areduce_nor_6_a2(
	.dataa(!fp_functions_0_areduce_nor_6_a0_combout),
	.datab(!fp_functions_0_areduce_nor_6_a1_combout),
	.datac(!fp_functions_0_areduce_nor_5_a0_combout),
	.datad(!fp_functions_0_arVStage_uid177_lzCountVal_uid85_fpAddTest_b_a0_a_a1_combout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_areduce_nor_6_a2_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_areduce_nor_6_a2.extended_lut = "off";
defparam fp_functions_0_areduce_nor_6_a2.lut_mask = 64'h0100010001000100;
defparam fp_functions_0_areduce_nor_6_a2.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_areduce_nor_6_a3(
	.dataa(!fp_functions_0_aredist1_vCount_uid152_lzCountVal_uid85_fpAddTest_q_1_q_a0_a_aq),
	.datab(!fp_functions_0_arVStage_uid165_lzCountVal_uid85_fpAddTest_merged_bit_select_b_a2_a_a4_combout),
	.datac(!fp_functions_0_arVStage_uid165_lzCountVal_uid85_fpAddTest_merged_bit_select_b_a3_a_a6_combout),
	.datad(!fp_functions_0_areduce_nor_6_a2_combout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_areduce_nor_6_a3_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_areduce_nor_6_a3.extended_lut = "off";
defparam fp_functions_0_areduce_nor_6_a3.lut_mask = 64'h0001000100010001;
defparam fp_functions_0_areduce_nor_6_a3.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_areduce_nor_8_a0(
	.dataa(!fp_functions_0_aredist18_exp_aSig_uid21_fpAddTest_b_2_q_a0_a_aq),
	.datab(!fp_functions_0_aredist18_exp_aSig_uid21_fpAddTest_b_2_q_a1_a_aq),
	.datac(!fp_functions_0_aredist18_exp_aSig_uid21_fpAddTest_b_2_q_a2_a_aq),
	.datad(!fp_functions_0_aredist18_exp_aSig_uid21_fpAddTest_b_2_q_a3_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_areduce_nor_8_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_areduce_nor_8_a0.extended_lut = "off";
defparam fp_functions_0_areduce_nor_8_a0.lut_mask = 64'h0001000100010001;
defparam fp_functions_0_areduce_nor_8_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_areduce_nor_8(
	.dataa(!fp_functions_0_aredist18_exp_aSig_uid21_fpAddTest_b_2_q_a4_a_aq),
	.datab(!fp_functions_0_aredist18_exp_aSig_uid21_fpAddTest_b_2_q_a5_a_aq),
	.datac(!fp_functions_0_aredist18_exp_aSig_uid21_fpAddTest_b_2_q_a6_a_aq),
	.datad(!fp_functions_0_aredist18_exp_aSig_uid21_fpAddTest_b_2_q_a7_a_aq),
	.datae(!fp_functions_0_areduce_nor_8_a0_combout),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_areduce_nor_8_acombout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_areduce_nor_8.extended_lut = "off";
defparam fp_functions_0_areduce_nor_8.lut_mask = 64'h0000000100000001;
defparam fp_functions_0_areduce_nor_8.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_areduce_nor_9_a0(
	.dataa(!fp_functions_0_aredist18_exp_aSig_uid21_fpAddTest_b_2_q_a0_a_aq),
	.datab(!fp_functions_0_aredist18_exp_aSig_uid21_fpAddTest_b_2_q_a1_a_aq),
	.datac(!fp_functions_0_aredist18_exp_aSig_uid21_fpAddTest_b_2_q_a2_a_aq),
	.datad(!fp_functions_0_aredist18_exp_aSig_uid21_fpAddTest_b_2_q_a3_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_areduce_nor_9_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_areduce_nor_9_a0.extended_lut = "off";
defparam fp_functions_0_areduce_nor_9_a0.lut_mask = 64'h8000800080008000;
defparam fp_functions_0_areduce_nor_9_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_areduce_nor_9(
	.dataa(!fp_functions_0_aredist18_exp_aSig_uid21_fpAddTest_b_2_q_a4_a_aq),
	.datab(!fp_functions_0_aredist18_exp_aSig_uid21_fpAddTest_b_2_q_a5_a_aq),
	.datac(!fp_functions_0_aredist18_exp_aSig_uid21_fpAddTest_b_2_q_a6_a_aq),
	.datad(!fp_functions_0_aredist18_exp_aSig_uid21_fpAddTest_b_2_q_a7_a_aq),
	.datae(!fp_functions_0_areduce_nor_9_a0_combout),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_areduce_nor_9_acombout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_areduce_nor_9.extended_lut = "off";
defparam fp_functions_0_areduce_nor_9.lut_mask = 64'h0000800000008000;
defparam fp_functions_0_areduce_nor_9.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aregInputs_uid118_fpAddTest_qi_a0_a_a1(
	.dataa(!fp_functions_0_aredist12_expXIsMax_uid38_fpAddTest_q_2_q_a0_a_aq),
	.datab(!fp_functions_0_aredist9_InvExpXIsZero_uid44_fpAddTest_q_2_q_a0_a_aq),
	.datac(!fp_functions_0_areduce_nor_8_acombout),
	.datad(!fp_functions_0_areduce_nor_9_acombout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aregInputs_uid118_fpAddTest_qi_a0_a_a1_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aregInputs_uid118_fpAddTest_qi_a0_a_a1.extended_lut = "off";
defparam fp_functions_0_aregInputs_uid118_fpAddTest_qi_a0_a_a1.lut_mask = 64'h2000200020002000;
defparam fp_functions_0_aregInputs_uid118_fpAddTest_qi_a0_a_a1.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aexcI_aSig_uid27_fpAddTest_q_a0_a(
	.dataa(!fp_functions_0_afracXIsZero_uid25_fpAddTest_delay_adelay_signals_a0_a_a0_a_aq),
	.datab(!fp_functions_0_areduce_nor_8_acombout),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aexcI_aSig_uid27_fpAddTest_q_a0_a_acombout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aexcI_aSig_uid27_fpAddTest_q_a0_a.extended_lut = "off";
defparam fp_functions_0_aexcI_aSig_uid27_fpAddTest_q_a0_a.lut_mask = 64'h1111111111111111;
defparam fp_functions_0_aexcI_aSig_uid27_fpAddTest_q_a0_a.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aexcI_bSig_uid41_fpAddTest_q_a0_a(
	.dataa(!fp_functions_0_aredist12_expXIsMax_uid38_fpAddTest_q_2_q_a0_a_aq),
	.datab(!fp_functions_0_aredist11_fracXIsZero_uid39_fpAddTest_q_2_q_a0_a_aq),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aexcI_bSig_uid41_fpAddTest_q_a0_a_acombout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aexcI_bSig_uid41_fpAddTest_q_a0_a.extended_lut = "off";
defparam fp_functions_0_aexcI_bSig_uid41_fpAddTest_q_a0_a.lut_mask = 64'h1111111111111111;
defparam fp_functions_0_aexcI_bSig_uid41_fpAddTest_q_a0_a.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aexcN_bSig_uid42_fpAddTest_qi_a0_a(
	.dataa(!fp_functions_0_aredist12_expXIsMax_uid38_fpAddTest_q_2_q_a0_a_aq),
	.datab(!fp_functions_0_aredist11_fracXIsZero_uid39_fpAddTest_q_2_q_a0_a_aq),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aexcN_bSig_uid42_fpAddTest_qi_a0_a_acombout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aexcN_bSig_uid42_fpAddTest_qi_a0_a.extended_lut = "off";
defparam fp_functions_0_aexcN_bSig_uid42_fpAddTest_qi_a0_a.lut_mask = 64'h4444444444444444;
defparam fp_functions_0_aexcN_bSig_uid42_fpAddTest_qi_a0_a.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aexcN_aSig_uid28_fpAddTest_qi_a0_a(
	.dataa(!fp_functions_0_afracXIsZero_uid25_fpAddTest_delay_adelay_signals_a0_a_a0_a_aq),
	.datab(!fp_functions_0_areduce_nor_8_acombout),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aexcN_aSig_uid28_fpAddTest_qi_a0_a_acombout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aexcN_aSig_uid28_fpAddTest_qi_a0_a.extended_lut = "off";
defparam fp_functions_0_aexcN_aSig_uid28_fpAddTest_qi_a0_a.lut_mask = 64'h2222222222222222;
defparam fp_functions_0_aexcN_aSig_uid28_fpAddTest_qi_a0_a.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_asignRInfRZRReg_uid137_fpAddTest_qi_a0_a_a1(
	.dataa(!fp_functions_0_afracXIsZero_uid25_fpAddTest_delay_adelay_signals_a0_a_a0_a_aq),
	.datab(!fp_functions_0_aredist13_excZ_bSig_uid17_uid37_fpAddTest_q_2_q_a0_a_aq),
	.datac(!fp_functions_0_aredist6_sigB_uid51_fpAddTest_b_2_q_a0_a_aq),
	.datad(!fp_functions_0_areduce_nor_8_acombout),
	.datae(!fp_functions_0_areduce_nor_9_acombout),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_asignRInfRZRReg_uid137_fpAddTest_qi_a0_a_a1_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_asignRInfRZRReg_uid137_fpAddTest_qi_a0_a_a1.extended_lut = "off";
defparam fp_functions_0_asignRInfRZRReg_uid137_fpAddTest_qi_a0_a_a1.lut_mask = 64'h3355035733550357;
defparam fp_functions_0_asignRInfRZRReg_uid137_fpAddTest_qi_a0_a_a1.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_asignRInfRZRReg_uid137_fpAddTest_qi_a0_a_a2(
	.dataa(!fp_functions_0_aredist6_sigB_uid51_fpAddTest_b_2_q_a0_a_aq),
	.datab(!fp_functions_0_aredist8_sigA_uid50_fpAddTest_b_2_q_a0_a_aq),
	.datac(!fp_functions_0_aexcI_bSig_uid41_fpAddTest_q_a0_a_acombout),
	.datad(!fp_functions_0_aregInputs_uid118_fpAddTest_qi_a0_a_a1_combout),
	.datae(!fp_functions_0_asignRInfRZRReg_uid137_fpAddTest_qi_a0_a_a1_combout),
	.dataf(!fp_functions_0_areduce_nor_6_a3_combout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_asignRInfRZRReg_uid137_fpAddTest_qi_a0_a_a2_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_asignRInfRZRReg_uid137_fpAddTest_qi_a0_a_a2.extended_lut = "off";
defparam fp_functions_0_asignRInfRZRReg_uid137_fpAddTest_qi_a0_a_a2.lut_mask = 64'h0537373705053737;
defparam fp_functions_0_asignRInfRZRReg_uid137_fpAddTest_qi_a0_a_a2.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai2460_a1(
	.dataa(!fp_functions_0_aadd_4_a11_sumout),
	.datab(!fp_functions_0_aadd_4_a16_sumout),
	.datac(!fp_functions_0_aadd_4_a21_sumout),
	.datad(!fp_functions_0_aadd_4_a26_sumout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai2460_a1_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai2460_a1.extended_lut = "off";
defparam fp_functions_0_ai2460_a1.lut_mask = 64'h8000800080008000;
defparam fp_functions_0_ai2460_a1.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai2460_a2(
	.dataa(!fp_functions_0_aadd_4_a6_sumout),
	.datab(!fp_functions_0_ai2460_a1_combout),
	.datac(!fp_functions_0_aadd_4_a31_sumout),
	.datad(!fp_functions_0_aadd_4_a36_sumout),
	.datae(!fp_functions_0_aadd_4_a41_sumout),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai2460_a2_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai2460_a2.extended_lut = "off";
defparam fp_functions_0_ai2460_a2.lut_mask = 64'h2000000020000000;
defparam fp_functions_0_ai2460_a2.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai2460_a3(
	.dataa(!fp_functions_0_aadd_4_a56_sumout),
	.datab(!fp_functions_0_aadd_4_a61_sumout),
	.datac(!fp_functions_0_aadd_4_a66_sumout),
	.datad(!fp_functions_0_aadd_4_a71_sumout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai2460_a3_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai2460_a3.extended_lut = "off";
defparam fp_functions_0_ai2460_a3.lut_mask = 64'h8000800080008000;
defparam fp_functions_0_ai2460_a3.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_areduce_nor_2(
	.dataa(!fp_functions_0_aadd_4_a1_sumout),
	.datab(!fp_functions_0_ai2460_a2_combout),
	.datac(!fp_functions_0_aadd_4_a46_sumout),
	.datad(!fp_functions_0_aadd_4_a51_sumout),
	.datae(!fp_functions_0_ai2460_a3_combout),
	.dataf(!fp_functions_0_aadd_4_a76_sumout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_areduce_nor_2_acombout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_areduce_nor_2.extended_lut = "off";
defparam fp_functions_0_areduce_nor_2.lut_mask = 64'h0000200000000000;
defparam fp_functions_0_areduce_nor_2.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai2460_a4(
	.dataa(!fp_functions_0_aadd_4_a56_sumout),
	.datab(!fp_functions_0_aadd_4_a61_sumout),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai2460_a4_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai2460_a4.extended_lut = "off";
defparam fp_functions_0_ai2460_a4.lut_mask = 64'h8888888888888888;
defparam fp_functions_0_ai2460_a4.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai2459_a1(
	.dataa(!fp_functions_0_aadd_4_a1_sumout),
	.datab(!fp_functions_0_aadd_4_a46_sumout),
	.datac(!fp_functions_0_aadd_4_a51_sumout),
	.datad(!fp_functions_0_aadd_4_a76_sumout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai2459_a1_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai2459_a1.extended_lut = "off";
defparam fp_functions_0_ai2459_a1.lut_mask = 64'h8000800080008000;
defparam fp_functions_0_ai2459_a1.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai2467_a0(
	.dataa(!fp_functions_0_aadd_4_a81_sumout),
	.datab(!fp_functions_0_ai2460_a2_combout),
	.datac(!fp_functions_0_ai2460_a4_combout),
	.datad(!fp_functions_0_aadd_4_a66_sumout),
	.datae(!fp_functions_0_aadd_4_a71_sumout),
	.dataf(!fp_functions_0_ai2459_a1_combout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai2467_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai2467_a0.extended_lut = "off";
defparam fp_functions_0_ai2467_a0.lut_mask = 64'h00FF00FF01FF00FF;
defparam fp_functions_0_ai2467_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai2460_a5(
	.dataa(!fp_functions_0_aadd_4_a66_sumout),
	.datab(!fp_functions_0_aadd_4_a71_sumout),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai2460_a5_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai2460_a5.extended_lut = "off";
defparam fp_functions_0_ai2460_a5.lut_mask = 64'h8888888888888888;
defparam fp_functions_0_ai2460_a5.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai2467_a1(
	.dataa(!fp_functions_0_aadd_4_a86_sumout),
	.datab(!fp_functions_0_aadd_4_a56_sumout),
	.datac(!fp_functions_0_aadd_4_a61_sumout),
	.datad(!fp_functions_0_ai2460_a2_combout),
	.datae(!fp_functions_0_ai2460_a5_combout),
	.dataf(!fp_functions_0_ai2459_a1_combout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai2467_a1_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai2467_a1.extended_lut = "off";
defparam fp_functions_0_ai2467_a1.lut_mask = 64'h0F0F0F0F0F0F0F4F;
defparam fp_functions_0_ai2467_a1.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai2460_a6(
	.dataa(!fp_functions_0_aadd_4_a46_sumout),
	.datab(!fp_functions_0_aadd_4_a51_sumout),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai2460_a6_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai2460_a6.extended_lut = "off";
defparam fp_functions_0_ai2460_a6.lut_mask = 64'h8888888888888888;
defparam fp_functions_0_ai2460_a6.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai2467_a2(
	.dataa(!fp_functions_0_aadd_4_a91_sumout),
	.datab(!fp_functions_0_aadd_4_a1_sumout),
	.datac(!fp_functions_0_ai2460_a2_combout),
	.datad(!fp_functions_0_ai2460_a3_combout),
	.datae(!fp_functions_0_ai2460_a6_combout),
	.dataf(!fp_functions_0_aadd_4_a76_sumout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai2467_a2_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai2467_a2.extended_lut = "off";
defparam fp_functions_0_ai2467_a2.lut_mask = 64'h3333333733333333;
defparam fp_functions_0_ai2467_a2.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai2467_a3(
	.dataa(!fp_functions_0_aadd_4_a96_sumout),
	.datab(!fp_functions_0_aadd_4_a56_sumout),
	.datac(!fp_functions_0_aadd_4_a61_sumout),
	.datad(!fp_functions_0_ai2460_a2_combout),
	.datae(!fp_functions_0_ai2460_a5_combout),
	.dataf(!fp_functions_0_ai2459_a1_combout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai2467_a3_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai2467_a3.extended_lut = "off";
defparam fp_functions_0_ai2467_a3.lut_mask = 64'h3333333333333373;
defparam fp_functions_0_ai2467_a3.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai2453_a1(
	.dataa(!fp_functions_0_aadd_4_a101_sumout),
	.datab(!fp_functions_0_aadd_4_a1_sumout),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai2453_a1_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai2453_a1.extended_lut = "off";
defparam fp_functions_0_ai2453_a1.lut_mask = 64'h4444444444444444;
defparam fp_functions_0_ai2453_a1.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai2467_a4(
	.dataa(!fp_functions_0_ai2453_a1_combout),
	.datab(!fp_functions_0_ai2460_a2_combout),
	.datac(!fp_functions_0_aadd_4_a46_sumout),
	.datad(!fp_functions_0_aadd_4_a51_sumout),
	.datae(!fp_functions_0_ai2460_a3_combout),
	.dataf(!fp_functions_0_aadd_4_a76_sumout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai2467_a4_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai2467_a4.extended_lut = "off";
defparam fp_functions_0_ai2467_a4.lut_mask = 64'h00001000FFFFFFFF;
defparam fp_functions_0_ai2467_a4.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai2454_a1(
	.dataa(!fp_functions_0_aadd_4_a106_sumout),
	.datab(!fp_functions_0_aadd_4_a46_sumout),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai2454_a1_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai2454_a1.extended_lut = "off";
defparam fp_functions_0_ai2454_a1.lut_mask = 64'h4444444444444444;
defparam fp_functions_0_ai2454_a1.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai2467_a5(
	.dataa(!fp_functions_0_aadd_4_a1_sumout),
	.datab(!fp_functions_0_ai2460_a2_combout),
	.datac(!fp_functions_0_aadd_4_a51_sumout),
	.datad(!fp_functions_0_ai2460_a3_combout),
	.datae(!fp_functions_0_ai2454_a1_combout),
	.dataf(!fp_functions_0_aadd_4_a76_sumout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai2467_a5_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai2467_a5.extended_lut = "off";
defparam fp_functions_0_ai2467_a5.lut_mask = 64'h0F0F0F2F0F0F0F0F;
defparam fp_functions_0_ai2467_a5.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai2460_a7(
	.dataa(!fp_functions_0_aadd_4_a6_sumout),
	.datab(!fp_functions_0_aadd_4_a31_sumout),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai2460_a7_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai2460_a7.extended_lut = "off";
defparam fp_functions_0_ai2460_a7.lut_mask = 64'h8888888888888888;
defparam fp_functions_0_ai2460_a7.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai2461_a1(
	.dataa(!fp_functions_0_aadd_4_a111_sumout),
	.datab(!fp_functions_0_aadd_4_a36_sumout),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai2461_a1_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai2461_a1.extended_lut = "off";
defparam fp_functions_0_ai2461_a1.lut_mask = 64'h4444444444444444;
defparam fp_functions_0_ai2461_a1.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai2467_a6(
	.dataa(!fp_functions_0_ai2460_a1_combout),
	.datab(!fp_functions_0_ai2460_a7_combout),
	.datac(!fp_functions_0_aadd_4_a41_sumout),
	.datad(!fp_functions_0_ai2461_a1_combout),
	.datae(!fp_functions_0_ai2460_a3_combout),
	.dataf(!fp_functions_0_ai2459_a1_combout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai2467_a6_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai2467_a6.extended_lut = "off";
defparam fp_functions_0_ai2467_a6.lut_mask = 64'h0F0F0F0F0F0F0F1F;
defparam fp_functions_0_ai2467_a6.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai2467_a7(
	.dataa(!fp_functions_0_aadd_4_a116_sumout),
	.datab(!fp_functions_0_ai2460_a2_combout),
	.datac(!fp_functions_0_ai2460_a4_combout),
	.datad(!fp_functions_0_aadd_4_a66_sumout),
	.datae(!fp_functions_0_aadd_4_a71_sumout),
	.dataf(!fp_functions_0_ai2459_a1_combout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai2467_a7_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai2467_a7.extended_lut = "off";
defparam fp_functions_0_ai2467_a7.lut_mask = 64'h0000FFFF0100FFFF;
defparam fp_functions_0_ai2467_a7.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai2455_a1(
	.dataa(!fp_functions_0_aadd_4_a121_sumout),
	.datab(!fp_functions_0_aadd_4_a51_sumout),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai2455_a1_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai2455_a1.extended_lut = "off";
defparam fp_functions_0_ai2455_a1.lut_mask = 64'h4444444444444444;
defparam fp_functions_0_ai2455_a1.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai2467_a8(
	.dataa(!fp_functions_0_aadd_4_a1_sumout),
	.datab(!fp_functions_0_ai2460_a2_combout),
	.datac(!fp_functions_0_aadd_4_a46_sumout),
	.datad(!fp_functions_0_ai2460_a3_combout),
	.datae(!fp_functions_0_aadd_4_a76_sumout),
	.dataf(!fp_functions_0_ai2455_a1_combout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai2467_a8_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai2467_a8.extended_lut = "off";
defparam fp_functions_0_ai2467_a8.lut_mask = 64'h0F0F0F0F0F2F0F0F;
defparam fp_functions_0_ai2467_a8.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai2462_a1(
	.dataa(!fp_functions_0_aadd_4_a126_sumout),
	.datab(!fp_functions_0_aadd_4_a41_sumout),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai2462_a1_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai2462_a1.extended_lut = "off";
defparam fp_functions_0_ai2462_a1.lut_mask = 64'h4444444444444444;
defparam fp_functions_0_ai2462_a1.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai2467_a9(
	.dataa(!fp_functions_0_ai2460_a1_combout),
	.datab(!fp_functions_0_ai2460_a7_combout),
	.datac(!fp_functions_0_aadd_4_a36_sumout),
	.datad(!fp_functions_0_ai2462_a1_combout),
	.datae(!fp_functions_0_ai2460_a3_combout),
	.dataf(!fp_functions_0_ai2459_a1_combout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai2467_a9_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai2467_a9.extended_lut = "off";
defparam fp_functions_0_ai2467_a9.lut_mask = 64'h0F0F0F0F0F0F0F1F;
defparam fp_functions_0_ai2467_a9.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai2463_a1(
	.dataa(!fp_functions_0_aadd_4_a131_sumout),
	.datab(!fp_functions_0_aadd_4_a6_sumout),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai2463_a1_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai2463_a1.extended_lut = "off";
defparam fp_functions_0_ai2463_a1.lut_mask = 64'h4444444444444444;
defparam fp_functions_0_ai2463_a1.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai2460_a8(
	.dataa(!fp_functions_0_aadd_4_a36_sumout),
	.datab(!fp_functions_0_aadd_4_a41_sumout),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai2460_a8_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai2460_a8.extended_lut = "off";
defparam fp_functions_0_ai2460_a8.lut_mask = 64'h8888888888888888;
defparam fp_functions_0_ai2460_a8.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai2467_a10(
	.dataa(!fp_functions_0_ai2460_a1_combout),
	.datab(!fp_functions_0_aadd_4_a31_sumout),
	.datac(!fp_functions_0_ai2463_a1_combout),
	.datad(!fp_functions_0_ai2460_a8_combout),
	.datae(!fp_functions_0_ai2460_a3_combout),
	.dataf(!fp_functions_0_ai2459_a1_combout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai2467_a10_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai2467_a10.extended_lut = "off";
defparam fp_functions_0_ai2467_a10.lut_mask = 64'h3333333333333337;
defparam fp_functions_0_ai2467_a10.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_areduce_nor_1_a0(
	.dataa(!fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a16_a_aq),
	.datab(!fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a0_a_aq),
	.datac(!fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a1_a_aq),
	.datad(!fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a9_a_aq),
	.datae(!fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a4_a_aq),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_areduce_nor_1_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_areduce_nor_1_a0.extended_lut = "off";
defparam fp_functions_0_areduce_nor_1_a0.lut_mask = 64'h8000000080000000;
defparam fp_functions_0_areduce_nor_1_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_areduce_nor_1_a1(
	.dataa(!fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a21_a_aq),
	.datab(!fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a20_a_aq),
	.datac(!fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a19_a_aq),
	.datad(!fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a17_a_aq),
	.datae(!fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a18_a_aq),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_areduce_nor_1_a1_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_areduce_nor_1_a1.extended_lut = "off";
defparam fp_functions_0_areduce_nor_1_a1.lut_mask = 64'h8000000080000000;
defparam fp_functions_0_areduce_nor_1_a1.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_areduce_nor_1_a2(
	.dataa(!fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a8_a_aq),
	.datab(!fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a7_a_aq),
	.datac(!fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a6_a_aq),
	.datad(!fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a5_a_aq),
	.datae(!fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a2_a_aq),
	.dataf(!fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a3_a_aq),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_areduce_nor_1_a2_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_areduce_nor_1_a2.extended_lut = "off";
defparam fp_functions_0_areduce_nor_1_a2.lut_mask = 64'h8000000000000000;
defparam fp_functions_0_areduce_nor_1_a2.shared_arith = "off";

fourteennm_ff fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a15_a(
	.clk(clk),
	.d(fp_functions_0_ai1783_a16_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a15_a_aq));
defparam fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a15_a.is_wysiwyg = "true";
defparam fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a15_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a14_a(
	.clk(clk),
	.d(fp_functions_0_ai1783_a17_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a14_a_aq));
defparam fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a14_a.is_wysiwyg = "true";
defparam fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a14_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a13_a(
	.clk(clk),
	.d(fp_functions_0_ai1783_a49_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a13_a_aq));
defparam fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a13_a.is_wysiwyg = "true";
defparam fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a13_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a12_a(
	.clk(clk),
	.d(fp_functions_0_ai1783_a44_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a12_a_aq));
defparam fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a12_a.is_wysiwyg = "true";
defparam fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a12_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a10_a(
	.clk(clk),
	.d(fp_functions_0_ai1783_a39_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a10_a_aq));
defparam fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a10_a.is_wysiwyg = "true";
defparam fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a10_a.power_up = "dont_care";

fourteennm_ff fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a11_a(
	.clk(clk),
	.d(fp_functions_0_ai1783_a34_combout),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.q(fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a11_a_aq));
defparam fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a11_a.is_wysiwyg = "true";
defparam fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a11_a.power_up = "dont_care";

fourteennm_lcell_comb fp_functions_0_areduce_nor_1_a3(
	.dataa(!fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a15_a_aq),
	.datab(!fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a14_a_aq),
	.datac(!fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a13_a_aq),
	.datad(!fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a12_a_aq),
	.datae(!fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a10_a_aq),
	.dataf(!fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a11_a_aq),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_areduce_nor_1_a3_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_areduce_nor_1_a3.extended_lut = "off";
defparam fp_functions_0_areduce_nor_1_a3.lut_mask = 64'h8000000000000000;
defparam fp_functions_0_areduce_nor_1_a3.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_areduce_nor_1_a4(
	.dataa(!fp_functions_0_ashiftedOut_uid63_fpAddTest_o_a10_a_aq),
	.datab(!fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a22_a_aq),
	.datac(!fp_functions_0_areduce_nor_1_a0_combout),
	.datad(!fp_functions_0_areduce_nor_1_a1_combout),
	.datae(!fp_functions_0_areduce_nor_1_a2_combout),
	.dataf(!fp_functions_0_areduce_nor_1_a3_combout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_areduce_nor_1_a4_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_areduce_nor_1_a4.extended_lut = "off";
defparam fp_functions_0_areduce_nor_1_a4.lut_mask = 64'hAAAAAAAAAAAAAAA2;
defparam fp_functions_0_areduce_nor_1_a4.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai2464_a1(
	.dataa(!fp_functions_0_areduce_nor_1_a4_combout),
	.datab(!fp_functions_0_aadd_4_a31_sumout),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai2464_a1_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai2464_a1.extended_lut = "off";
defparam fp_functions_0_ai2464_a1.lut_mask = 64'h4444444444444444;
defparam fp_functions_0_ai2464_a1.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai2467_a11(
	.dataa(!fp_functions_0_aadd_4_a6_sumout),
	.datab(!fp_functions_0_ai2460_a1_combout),
	.datac(!fp_functions_0_ai2464_a1_combout),
	.datad(!fp_functions_0_ai2460_a8_combout),
	.datae(!fp_functions_0_ai2460_a3_combout),
	.dataf(!fp_functions_0_ai2459_a1_combout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai2467_a11_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai2467_a11.extended_lut = "off";
defparam fp_functions_0_ai2467_a11.lut_mask = 64'h5555555555555557;
defparam fp_functions_0_ai2467_a11.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai2460_a9(
	.dataa(!fp_functions_0_aadd_4_a11_sumout),
	.datab(!fp_functions_0_aadd_4_a16_sumout),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai2460_a9_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai2460_a9.extended_lut = "off";
defparam fp_functions_0_ai2460_a9.lut_mask = 64'h8888888888888888;
defparam fp_functions_0_ai2460_a9.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai2460_a10(
	.dataa(!fp_functions_0_aadd_4_a6_sumout),
	.datab(!fp_functions_0_aadd_4_a31_sumout),
	.datac(!fp_functions_0_aadd_4_a36_sumout),
	.datad(!fp_functions_0_aadd_4_a41_sumout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai2460_a10_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai2460_a10.extended_lut = "off";
defparam fp_functions_0_ai2460_a10.lut_mask = 64'h8000800080008000;
defparam fp_functions_0_ai2460_a10.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai2467_a12(
	.dataa(!fp_functions_0_ai2460_a9_combout),
	.datab(!fp_functions_0_aadd_4_a21_sumout),
	.datac(!fp_functions_0_aadd_4_a26_sumout),
	.datad(!fp_functions_0_ai2460_a10_combout),
	.datae(!fp_functions_0_ai2460_a3_combout),
	.dataf(!fp_functions_0_ai2459_a1_combout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai2467_a12_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai2467_a12.extended_lut = "off";
defparam fp_functions_0_ai2467_a12.lut_mask = 64'h0F0F0F0F0F0F0F4F;
defparam fp_functions_0_ai2467_a12.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai2467_a13(
	.dataa(!fp_functions_0_ai2460_a9_combout),
	.datab(!fp_functions_0_aadd_4_a21_sumout),
	.datac(!fp_functions_0_aadd_4_a26_sumout),
	.datad(!fp_functions_0_ai2460_a10_combout),
	.datae(!fp_functions_0_ai2460_a3_combout),
	.dataf(!fp_functions_0_ai2459_a1_combout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai2467_a13_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai2467_a13.extended_lut = "off";
defparam fp_functions_0_ai2467_a13.lut_mask = 64'h3333333333333373;
defparam fp_functions_0_ai2467_a13.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai2467_a14(
	.dataa(!fp_functions_0_aadd_4_a11_sumout),
	.datab(!fp_functions_0_aadd_4_a21_sumout),
	.datac(!fp_functions_0_aadd_4_a26_sumout),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai2467_a14_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai2467_a14.extended_lut = "off";
defparam fp_functions_0_ai2467_a14.lut_mask = 64'h8080808080808080;
defparam fp_functions_0_ai2467_a14.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai2467_a15(
	.dataa(!fp_functions_0_aadd_4_a16_sumout),
	.datab(!fp_functions_0_ai2467_a14_combout),
	.datac(!fp_functions_0_ai2460_a10_combout),
	.datad(!fp_functions_0_ai2460_a3_combout),
	.datae(!fp_functions_0_ai2459_a1_combout),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai2467_a15_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai2467_a15.extended_lut = "off";
defparam fp_functions_0_ai2467_a15.lut_mask = 64'h5555555755555557;
defparam fp_functions_0_ai2467_a15.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_afracBAddOpPostXor_uid81_fpAddTest_b_a26_a(
	.dataa(!fp_functions_0_aredist7_sigA_uid50_fpAddTest_b_1_q_a0_a_aq),
	.datab(!fp_functions_0_aredist5_sigB_uid51_fpAddTest_b_1_q_a0_a_aq),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_afracBAddOpPostXor_uid81_fpAddTest_b_a26_a_acombout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_afracBAddOpPostXor_uid81_fpAddTest_b_a26_a.extended_lut = "off";
defparam fp_functions_0_afracBAddOpPostXor_uid81_fpAddTest_b_a26_a.lut_mask = 64'h6666666666666666;
defparam fp_functions_0_afracBAddOpPostXor_uid81_fpAddTest_b_a26_a.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_areduce_nor_11_a0(
	.dataa(!fp_functions_0_aredist17_frac_aSig_uid22_fpAddTest_b_1_q_a15_a_aq),
	.datab(!fp_functions_0_aredist17_frac_aSig_uid22_fpAddTest_b_1_q_a16_a_aq),
	.datac(!fp_functions_0_aredist17_frac_aSig_uid22_fpAddTest_b_1_q_a17_a_aq),
	.datad(!fp_functions_0_aredist17_frac_aSig_uid22_fpAddTest_b_1_q_a18_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_areduce_nor_11_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_areduce_nor_11_a0.extended_lut = "off";
defparam fp_functions_0_areduce_nor_11_a0.lut_mask = 64'h8000800080008000;
defparam fp_functions_0_areduce_nor_11_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_areduce_nor_11_a1(
	.dataa(!fp_functions_0_aredist17_frac_aSig_uid22_fpAddTest_b_1_q_a20_a_aq),
	.datab(!fp_functions_0_aredist17_frac_aSig_uid22_fpAddTest_b_1_q_a22_a_aq),
	.datac(!fp_functions_0_aredist17_frac_aSig_uid22_fpAddTest_b_1_q_a2_a_aq),
	.datad(!fp_functions_0_aredist17_frac_aSig_uid22_fpAddTest_b_1_q_a0_a_aq),
	.datae(!fp_functions_0_aredist17_frac_aSig_uid22_fpAddTest_b_1_q_a1_a_aq),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_areduce_nor_11_a1_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_areduce_nor_11_a1.extended_lut = "off";
defparam fp_functions_0_areduce_nor_11_a1.lut_mask = 64'h8000000080000000;
defparam fp_functions_0_areduce_nor_11_a1.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_areduce_nor_11_a2(
	.dataa(!fp_functions_0_aredist17_frac_aSig_uid22_fpAddTest_b_1_q_a9_a_aq),
	.datab(!fp_functions_0_aredist17_frac_aSig_uid22_fpAddTest_b_1_q_a10_a_aq),
	.datac(!fp_functions_0_aredist17_frac_aSig_uid22_fpAddTest_b_1_q_a11_a_aq),
	.datad(!fp_functions_0_aredist17_frac_aSig_uid22_fpAddTest_b_1_q_a12_a_aq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_areduce_nor_11_a2_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_areduce_nor_11_a2.extended_lut = "off";
defparam fp_functions_0_areduce_nor_11_a2.lut_mask = 64'h8000800080008000;
defparam fp_functions_0_areduce_nor_11_a2.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_areduce_nor_11_a3(
	.dataa(!fp_functions_0_aredist17_frac_aSig_uid22_fpAddTest_b_1_q_a3_a_aq),
	.datab(!fp_functions_0_aredist17_frac_aSig_uid22_fpAddTest_b_1_q_a4_a_aq),
	.datac(!fp_functions_0_aredist17_frac_aSig_uid22_fpAddTest_b_1_q_a5_a_aq),
	.datad(!fp_functions_0_aredist17_frac_aSig_uid22_fpAddTest_b_1_q_a6_a_aq),
	.datae(!fp_functions_0_aredist17_frac_aSig_uid22_fpAddTest_b_1_q_a7_a_aq),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_areduce_nor_11_a3_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_areduce_nor_11_a3.extended_lut = "off";
defparam fp_functions_0_areduce_nor_11_a3.lut_mask = 64'h8000000080000000;
defparam fp_functions_0_areduce_nor_11_a3.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_areduce_nor_11_a4(
	.dataa(!fp_functions_0_aredist17_frac_aSig_uid22_fpAddTest_b_1_q_a8_a_aq),
	.datab(!fp_functions_0_aredist17_frac_aSig_uid22_fpAddTest_b_1_q_a13_a_aq),
	.datac(!fp_functions_0_aredist17_frac_aSig_uid22_fpAddTest_b_1_q_a14_a_aq),
	.datad(!fp_functions_0_areduce_nor_11_a2_combout),
	.datae(!fp_functions_0_areduce_nor_11_a3_combout),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_areduce_nor_11_a4_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_areduce_nor_11_a4.extended_lut = "off";
defparam fp_functions_0_areduce_nor_11_a4.lut_mask = 64'h0000008000000080;
defparam fp_functions_0_areduce_nor_11_a4.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_areduce_nor_11(
	.dataa(!fp_functions_0_aredist17_frac_aSig_uid22_fpAddTest_b_1_q_a19_a_aq),
	.datab(!fp_functions_0_aredist17_frac_aSig_uid22_fpAddTest_b_1_q_a21_a_aq),
	.datac(!fp_functions_0_areduce_nor_11_a0_combout),
	.datad(!fp_functions_0_areduce_nor_11_a1_combout),
	.datae(!fp_functions_0_areduce_nor_11_a4_combout),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_areduce_nor_11_acombout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_areduce_nor_11.extended_lut = "off";
defparam fp_functions_0_areduce_nor_11.lut_mask = 64'h0000000800000008;
defparam fp_functions_0_areduce_nor_11.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_areduce_nor_4(
	.dataa(!fp_functions_0_areduce_nor_6_a0_combout),
	.datab(!fp_functions_0_arVStage_uid165_lzCountVal_uid85_fpAddTest_merged_bit_select_b_a3_a_a6_combout),
	.datac(!fp_functions_0_areduce_nor_6_a1_combout),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_areduce_nor_4_acombout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_areduce_nor_4.extended_lut = "off";
defparam fp_functions_0_areduce_nor_4.lut_mask = 64'hFEFEFEFEFEFEFEFE;
defparam fp_functions_0_areduce_nor_4.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_areduce_nor_3(
	.dataa(!fp_functions_0_avStagei_uid157_lzCountVal_uid85_fpAddTest_q_a15_a_aq),
	.datab(!fp_functions_0_avStagei_uid157_lzCountVal_uid85_fpAddTest_q_a14_a_aq),
	.datac(!fp_functions_0_arVStage_uid165_lzCountVal_uid85_fpAddTest_merged_bit_select_b_a2_a_a5_combout),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_areduce_nor_3_acombout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_areduce_nor_3.extended_lut = "off";
defparam fp_functions_0_areduce_nor_3.lut_mask = 64'hF7F7F7F7F7F7F7F7;
defparam fp_functions_0_areduce_nor_3.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_186_a0(
	.dataa(!fp_functions_0_aredist1_vCount_uid152_lzCountVal_uid85_fpAddTest_q_1_q_a0_a_aq),
	.datab(!fp_functions_0_aredist0_vStage_uid154_lzCountVal_uid85_fpAddTest_b_1_q_a0_a_aq),
	.datac(!fp_functions_0_areduce_nor_3_acombout),
	.datad(!fp_functions_0_areduce_nor_5_a0_combout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_186_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_186_a0.extended_lut = "off";
defparam fp_functions_0_aMux_186_a0.lut_mask = 64'h0002000200020002;
defparam fp_functions_0_aMux_186_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_186_a1(
	.dataa(!fp_functions_0_aredist1_vCount_uid152_lzCountVal_uid85_fpAddTest_q_1_q_a0_a_aq),
	.datab(!fp_functions_0_aredist0_vStage_uid154_lzCountVal_uid85_fpAddTest_b_1_q_a3_a_aq),
	.datac(!fp_functions_0_aredist0_vStage_uid154_lzCountVal_uid85_fpAddTest_b_1_q_a1_a_aq),
	.datad(!fp_functions_0_areduce_nor_3_acombout),
	.datae(!fp_functions_0_areduce_nor_5_a0_combout),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_186_a1_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_186_a1.extended_lut = "off";
defparam fp_functions_0_aMux_186_a1.lut_mask = 64'h000A0022000A0022;
defparam fp_functions_0_aMux_186_a1.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_186_a2(
	.dataa(!fp_functions_0_aredist1_vCount_uid152_lzCountVal_uid85_fpAddTest_q_1_q_a0_a_aq),
	.datab(!fp_functions_0_aredist0_vStage_uid154_lzCountVal_uid85_fpAddTest_b_1_q_a4_a_aq),
	.datac(!fp_functions_0_aredist0_vStage_uid154_lzCountVal_uid85_fpAddTest_b_1_q_a2_a_aq),
	.datad(!fp_functions_0_areduce_nor_3_acombout),
	.datae(!fp_functions_0_areduce_nor_5_a0_combout),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_186_a2_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_186_a2.extended_lut = "off";
defparam fp_functions_0_aMux_186_a2.lut_mask = 64'h000A0022000A0022;
defparam fp_functions_0_aMux_186_a2.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai3337_a0(
	.dataa(!fp_functions_0_areduce_nor_4_acombout),
	.datab(!fp_functions_0_arVStage_uid177_lzCountVal_uid85_fpAddTest_b_a0_a_a1_combout),
	.datac(!fp_functions_0_aMux_186_a0_combout),
	.datad(!fp_functions_0_aMux_186_a1_combout),
	.datae(!fp_functions_0_aMux_186_a2_combout),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai3337_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai3337_a0.extended_lut = "off";
defparam fp_functions_0_ai3337_a0.lut_mask = 64'h08194C5D08194C5D;
defparam fp_functions_0_ai3337_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_areduce_nor_12(
	.dataa(!fp_functions_0_aleftShiftStage2_uid249_fracPostNormExt_uid88_fpAddTest_q_a4_a_aq),
	.datab(!fp_functions_0_aleftShiftStage2_uid249_fracPostNormExt_uid88_fpAddTest_q_a3_a_aq),
	.datac(!fp_functions_0_aleftShiftStage2_uid249_fracPostNormExt_uid88_fpAddTest_q_a2_a_aq),
	.datad(!fp_functions_0_aleftShiftStage2_uid249_fracPostNormExt_uid88_fpAddTest_q_a0_a_aq),
	.datae(!fp_functions_0_aleftShiftStage2_uid249_fracPostNormExt_uid88_fpAddTest_q_a1_a_aq),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_areduce_nor_12_acombout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_areduce_nor_12.extended_lut = "off";
defparam fp_functions_0_areduce_nor_12.lut_mask = 64'hDFFFFFFFDFFFFFFF;
defparam fp_functions_0_areduce_nor_12.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_186_a3(
	.dataa(!fp_functions_0_aredist1_vCount_uid152_lzCountVal_uid85_fpAddTest_q_1_q_a0_a_aq),
	.datab(!fp_functions_0_aredist0_vStage_uid154_lzCountVal_uid85_fpAddTest_b_1_q_a1_a_aq),
	.datac(!fp_functions_0_areduce_nor_3_acombout),
	.datad(!fp_functions_0_areduce_nor_5_a0_combout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_186_a3_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_186_a3.extended_lut = "off";
defparam fp_functions_0_aMux_186_a3.lut_mask = 64'h0002000200020002;
defparam fp_functions_0_aMux_186_a3.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_186_a4(
	.dataa(!fp_functions_0_aredist1_vCount_uid152_lzCountVal_uid85_fpAddTest_q_1_q_a0_a_aq),
	.datab(!fp_functions_0_aredist0_vStage_uid154_lzCountVal_uid85_fpAddTest_b_1_q_a3_a_aq),
	.datac(!fp_functions_0_aredist0_vStage_uid154_lzCountVal_uid85_fpAddTest_b_1_q_a5_a_aq),
	.datad(!fp_functions_0_areduce_nor_3_acombout),
	.datae(!fp_functions_0_areduce_nor_5_a0_combout),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_186_a4_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_186_a4.extended_lut = "off";
defparam fp_functions_0_aMux_186_a4.lut_mask = 64'h0022000A0022000A;
defparam fp_functions_0_aMux_186_a4.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai3365_a0(
	.dataa(!fp_functions_0_aMux_186_a0_combout),
	.datab(!fp_functions_0_aMux_186_a2_combout),
	.datac(!fp_functions_0_aMux_186_a3_combout),
	.datad(!fp_functions_0_aMux_186_a4_combout),
	.datae(!fp_functions_0_areduce_nor_4_acombout),
	.dataf(!fp_functions_0_arVStage_uid177_lzCountVal_uid85_fpAddTest_b_a0_a_a1_combout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai3365_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai3365_a0.extended_lut = "off";
defparam fp_functions_0_ai3365_a0.lut_mask = 64'h0F0F00FF55553333;
defparam fp_functions_0_ai3365_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_186_a5(
	.dataa(!fp_functions_0_aredist1_vCount_uid152_lzCountVal_uid85_fpAddTest_q_1_q_a0_a_aq),
	.datab(!fp_functions_0_aredist0_vStage_uid154_lzCountVal_uid85_fpAddTest_b_1_q_a0_a_aq),
	.datac(!fp_functions_0_aredist0_vStage_uid154_lzCountVal_uid85_fpAddTest_b_1_q_a2_a_aq),
	.datad(!fp_functions_0_areduce_nor_3_acombout),
	.datae(!fp_functions_0_areduce_nor_5_a0_combout),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_186_a5_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_186_a5.extended_lut = "off";
defparam fp_functions_0_aMux_186_a5.lut_mask = 64'h0022000A0022000A;
defparam fp_functions_0_aMux_186_a5.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_186_a6(
	.dataa(!fp_functions_0_aredist1_vCount_uid152_lzCountVal_uid85_fpAddTest_q_1_q_a0_a_aq),
	.datab(!fp_functions_0_aredist0_vStage_uid154_lzCountVal_uid85_fpAddTest_b_1_q_a4_a_aq),
	.datac(!fp_functions_0_aredist0_vStage_uid154_lzCountVal_uid85_fpAddTest_b_1_q_a6_a_aq),
	.datad(!fp_functions_0_areduce_nor_3_acombout),
	.datae(!fp_functions_0_areduce_nor_5_a0_combout),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_186_a6_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_186_a6.extended_lut = "off";
defparam fp_functions_0_aMux_186_a6.lut_mask = 64'h0022000A0022000A;
defparam fp_functions_0_aMux_186_a6.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai3365_a1(
	.dataa(!fp_functions_0_aMux_186_a3_combout),
	.datab(!fp_functions_0_aMux_186_a4_combout),
	.datac(!fp_functions_0_aMux_186_a5_combout),
	.datad(!fp_functions_0_aMux_186_a6_combout),
	.datae(!fp_functions_0_areduce_nor_4_acombout),
	.dataf(!fp_functions_0_arVStage_uid177_lzCountVal_uid85_fpAddTest_b_a0_a_a1_combout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai3365_a1_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai3365_a1.extended_lut = "off";
defparam fp_functions_0_ai3365_a1.lut_mask = 64'h0F0F00FF55553333;
defparam fp_functions_0_ai3365_a1.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_186_a7(
	.dataa(!fp_functions_0_aredist1_vCount_uid152_lzCountVal_uid85_fpAddTest_q_1_q_a0_a_aq),
	.datab(!fp_functions_0_aredist0_vStage_uid154_lzCountVal_uid85_fpAddTest_b_1_q_a5_a_aq),
	.datac(!fp_functions_0_aredist0_vStage_uid154_lzCountVal_uid85_fpAddTest_b_1_q_a7_a_aq),
	.datad(!fp_functions_0_areduce_nor_3_acombout),
	.datae(!fp_functions_0_areduce_nor_5_a0_combout),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_186_a7_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_186_a7.extended_lut = "off";
defparam fp_functions_0_aMux_186_a7.lut_mask = 64'h0022000A0022000A;
defparam fp_functions_0_aMux_186_a7.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai3365_a2(
	.dataa(!fp_functions_0_aMux_186_a5_combout),
	.datab(!fp_functions_0_aMux_186_a6_combout),
	.datac(!fp_functions_0_aMux_186_a1_combout),
	.datad(!fp_functions_0_aMux_186_a7_combout),
	.datae(!fp_functions_0_areduce_nor_4_acombout),
	.dataf(!fp_functions_0_arVStage_uid177_lzCountVal_uid85_fpAddTest_b_a0_a_a1_combout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai3365_a2_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai3365_a2.extended_lut = "off";
defparam fp_functions_0_ai3365_a2.lut_mask = 64'h0F0F00FF55553333;
defparam fp_functions_0_ai3365_a2.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_186_a8(
	.dataa(!fp_functions_0_aredist0_vStage_uid154_lzCountVal_uid85_fpAddTest_b_1_q_a0_a_aq),
	.datab(!fp_functions_0_aredist0_vStage_uid154_lzCountVal_uid85_fpAddTest_b_1_q_a8_a_aq),
	.datac(!fp_functions_0_areduce_nor_3_acombout),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_186_a8_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_186_a8.extended_lut = "off";
defparam fp_functions_0_aMux_186_a8.lut_mask = 64'h5353535353535353;
defparam fp_functions_0_aMux_186_a8.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_186_a9(
	.dataa(!fp_functions_0_aredist1_vCount_uid152_lzCountVal_uid85_fpAddTest_q_1_q_a0_a_aq),
	.datab(!fp_functions_0_aredist0_vStage_uid154_lzCountVal_uid85_fpAddTest_b_1_q_a6_a_aq),
	.datac(!fp_functions_0_areduce_nor_3_acombout),
	.datad(!fp_functions_0_aMux_186_a8_combout),
	.datae(!fp_functions_0_areduce_nor_5_a0_combout),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_186_a9_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_186_a9.extended_lut = "off";
defparam fp_functions_0_aMux_186_a9.lut_mask = 64'h020200AA020200AA;
defparam fp_functions_0_aMux_186_a9.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai3365_a3(
	.dataa(!fp_functions_0_aMux_186_a1_combout),
	.datab(!fp_functions_0_aMux_186_a7_combout),
	.datac(!fp_functions_0_aMux_186_a2_combout),
	.datad(!fp_functions_0_aMux_186_a9_combout),
	.datae(!fp_functions_0_areduce_nor_4_acombout),
	.dataf(!fp_functions_0_arVStage_uid177_lzCountVal_uid85_fpAddTest_b_a0_a_a1_combout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai3365_a3_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai3365_a3.extended_lut = "off";
defparam fp_functions_0_ai3365_a3.lut_mask = 64'h0F0F00FF55553333;
defparam fp_functions_0_ai3365_a3.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_186_a10(
	.dataa(!fp_functions_0_aredist0_vStage_uid154_lzCountVal_uid85_fpAddTest_b_1_q_a1_a_aq),
	.datab(!fp_functions_0_aredist0_vStage_uid154_lzCountVal_uid85_fpAddTest_b_1_q_a9_a_aq),
	.datac(!fp_functions_0_areduce_nor_3_acombout),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_186_a10_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_186_a10.extended_lut = "off";
defparam fp_functions_0_aMux_186_a10.lut_mask = 64'h5353535353535353;
defparam fp_functions_0_aMux_186_a10.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_186_a11(
	.dataa(!fp_functions_0_aredist1_vCount_uid152_lzCountVal_uid85_fpAddTest_q_1_q_a0_a_aq),
	.datab(!fp_functions_0_aredist0_vStage_uid154_lzCountVal_uid85_fpAddTest_b_1_q_a7_a_aq),
	.datac(!fp_functions_0_areduce_nor_3_acombout),
	.datad(!fp_functions_0_aMux_186_a10_combout),
	.datae(!fp_functions_0_areduce_nor_5_a0_combout),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_186_a11_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_186_a11.extended_lut = "off";
defparam fp_functions_0_aMux_186_a11.lut_mask = 64'h020200AA020200AA;
defparam fp_functions_0_aMux_186_a11.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai3365_a4(
	.dataa(!fp_functions_0_aMux_186_a2_combout),
	.datab(!fp_functions_0_aMux_186_a9_combout),
	.datac(!fp_functions_0_aMux_186_a4_combout),
	.datad(!fp_functions_0_aMux_186_a11_combout),
	.datae(!fp_functions_0_areduce_nor_4_acombout),
	.dataf(!fp_functions_0_arVStage_uid177_lzCountVal_uid85_fpAddTest_b_a0_a_a1_combout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai3365_a4_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai3365_a4.extended_lut = "off";
defparam fp_functions_0_ai3365_a4.lut_mask = 64'h0F0F00FF55553333;
defparam fp_functions_0_ai3365_a4.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_186_a12(
	.dataa(!fp_functions_0_aredist0_vStage_uid154_lzCountVal_uid85_fpAddTest_b_1_q_a2_a_aq),
	.datab(!fp_functions_0_aredist0_vStage_uid154_lzCountVal_uid85_fpAddTest_b_1_q_a10_a_aq),
	.datac(!fp_functions_0_areduce_nor_3_acombout),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_186_a12_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_186_a12.extended_lut = "off";
defparam fp_functions_0_aMux_186_a12.lut_mask = 64'h5353535353535353;
defparam fp_functions_0_aMux_186_a12.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_186_a13(
	.dataa(!fp_functions_0_aredist1_vCount_uid152_lzCountVal_uid85_fpAddTest_q_1_q_a0_a_aq),
	.datab(!fp_functions_0_aMux_186_a8_combout),
	.datac(!fp_functions_0_aMux_186_a12_combout),
	.datad(!fp_functions_0_areduce_nor_5_a0_combout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_186_a13_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_186_a13.extended_lut = "off";
defparam fp_functions_0_aMux_186_a13.lut_mask = 64'h220A220A220A220A;
defparam fp_functions_0_aMux_186_a13.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai3365_a5(
	.dataa(!fp_functions_0_aMux_186_a4_combout),
	.datab(!fp_functions_0_aMux_186_a11_combout),
	.datac(!fp_functions_0_aMux_186_a6_combout),
	.datad(!fp_functions_0_aMux_186_a13_combout),
	.datae(!fp_functions_0_areduce_nor_4_acombout),
	.dataf(!fp_functions_0_arVStage_uid177_lzCountVal_uid85_fpAddTest_b_a0_a_a1_combout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai3365_a5_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai3365_a5.extended_lut = "off";
defparam fp_functions_0_ai3365_a5.lut_mask = 64'h0F0F00FF55553333;
defparam fp_functions_0_ai3365_a5.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_186_a14(
	.dataa(!fp_functions_0_aredist0_vStage_uid154_lzCountVal_uid85_fpAddTest_b_1_q_a3_a_aq),
	.datab(!fp_functions_0_aredist3_fracGRS_uid84_fpAddTest_q_1_q_a11_a_aq),
	.datac(!fp_functions_0_areduce_nor_3_acombout),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_186_a14_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_186_a14.extended_lut = "off";
defparam fp_functions_0_aMux_186_a14.lut_mask = 64'h5353535353535353;
defparam fp_functions_0_aMux_186_a14.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_186_a15(
	.dataa(!fp_functions_0_aredist1_vCount_uid152_lzCountVal_uid85_fpAddTest_q_1_q_a0_a_aq),
	.datab(!fp_functions_0_aMux_186_a10_combout),
	.datac(!fp_functions_0_aMux_186_a14_combout),
	.datad(!fp_functions_0_areduce_nor_5_a0_combout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_186_a15_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_186_a15.extended_lut = "off";
defparam fp_functions_0_aMux_186_a15.lut_mask = 64'h220A220A220A220A;
defparam fp_functions_0_aMux_186_a15.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai3365_a6(
	.dataa(!fp_functions_0_aMux_186_a6_combout),
	.datab(!fp_functions_0_aMux_186_a13_combout),
	.datac(!fp_functions_0_aMux_186_a7_combout),
	.datad(!fp_functions_0_aMux_186_a15_combout),
	.datae(!fp_functions_0_areduce_nor_4_acombout),
	.dataf(!fp_functions_0_arVStage_uid177_lzCountVal_uid85_fpAddTest_b_a0_a_a1_combout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai3365_a6_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai3365_a6.extended_lut = "off";
defparam fp_functions_0_ai3365_a6.lut_mask = 64'h0F0F00FF55553333;
defparam fp_functions_0_ai3365_a6.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_186_a16(
	.dataa(!fp_functions_0_aredist0_vStage_uid154_lzCountVal_uid85_fpAddTest_b_1_q_a4_a_aq),
	.datab(!fp_functions_0_aredist3_fracGRS_uid84_fpAddTest_q_1_q_a12_a_aq),
	.datac(!fp_functions_0_areduce_nor_3_acombout),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_186_a16_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_186_a16.extended_lut = "off";
defparam fp_functions_0_aMux_186_a16.lut_mask = 64'h5353535353535353;
defparam fp_functions_0_aMux_186_a16.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_186_a17(
	.dataa(!fp_functions_0_aredist1_vCount_uid152_lzCountVal_uid85_fpAddTest_q_1_q_a0_a_aq),
	.datab(!fp_functions_0_aMux_186_a12_combout),
	.datac(!fp_functions_0_aMux_186_a16_combout),
	.datad(!fp_functions_0_areduce_nor_5_a0_combout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_186_a17_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_186_a17.extended_lut = "off";
defparam fp_functions_0_aMux_186_a17.lut_mask = 64'h220A220A220A220A;
defparam fp_functions_0_aMux_186_a17.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai3365_a7(
	.dataa(!fp_functions_0_aMux_186_a7_combout),
	.datab(!fp_functions_0_aMux_186_a15_combout),
	.datac(!fp_functions_0_aMux_186_a9_combout),
	.datad(!fp_functions_0_aMux_186_a17_combout),
	.datae(!fp_functions_0_areduce_nor_4_acombout),
	.dataf(!fp_functions_0_arVStage_uid177_lzCountVal_uid85_fpAddTest_b_a0_a_a1_combout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai3365_a7_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai3365_a7.extended_lut = "off";
defparam fp_functions_0_ai3365_a7.lut_mask = 64'h0F0F00FF55553333;
defparam fp_functions_0_ai3365_a7.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_186_a18(
	.dataa(!fp_functions_0_aredist0_vStage_uid154_lzCountVal_uid85_fpAddTest_b_1_q_a5_a_aq),
	.datab(!fp_functions_0_aredist3_fracGRS_uid84_fpAddTest_q_1_q_a13_a_aq),
	.datac(!fp_functions_0_areduce_nor_3_acombout),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_186_a18_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_186_a18.extended_lut = "off";
defparam fp_functions_0_aMux_186_a18.lut_mask = 64'h5353535353535353;
defparam fp_functions_0_aMux_186_a18.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_186_a19(
	.dataa(!fp_functions_0_aredist1_vCount_uid152_lzCountVal_uid85_fpAddTest_q_1_q_a0_a_aq),
	.datab(!fp_functions_0_aMux_186_a14_combout),
	.datac(!fp_functions_0_aMux_186_a18_combout),
	.datad(!fp_functions_0_areduce_nor_5_a0_combout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_186_a19_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_186_a19.extended_lut = "off";
defparam fp_functions_0_aMux_186_a19.lut_mask = 64'h220A220A220A220A;
defparam fp_functions_0_aMux_186_a19.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai3365_a8(
	.dataa(!fp_functions_0_aMux_186_a9_combout),
	.datab(!fp_functions_0_aMux_186_a17_combout),
	.datac(!fp_functions_0_aMux_186_a11_combout),
	.datad(!fp_functions_0_aMux_186_a19_combout),
	.datae(!fp_functions_0_areduce_nor_4_acombout),
	.dataf(!fp_functions_0_arVStage_uid177_lzCountVal_uid85_fpAddTest_b_a0_a_a1_combout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai3365_a8_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai3365_a8.extended_lut = "off";
defparam fp_functions_0_ai3365_a8.lut_mask = 64'h0F0F00FF55553333;
defparam fp_functions_0_ai3365_a8.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_186_a20(
	.dataa(!fp_functions_0_aredist0_vStage_uid154_lzCountVal_uid85_fpAddTest_b_1_q_a6_a_aq),
	.datab(!fp_functions_0_aredist3_fracGRS_uid84_fpAddTest_q_1_q_a14_a_aq),
	.datac(!fp_functions_0_areduce_nor_3_acombout),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_186_a20_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_186_a20.extended_lut = "off";
defparam fp_functions_0_aMux_186_a20.lut_mask = 64'h5353535353535353;
defparam fp_functions_0_aMux_186_a20.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_186_a21(
	.dataa(!fp_functions_0_aredist1_vCount_uid152_lzCountVal_uid85_fpAddTest_q_1_q_a0_a_aq),
	.datab(!fp_functions_0_aMux_186_a16_combout),
	.datac(!fp_functions_0_aMux_186_a20_combout),
	.datad(!fp_functions_0_areduce_nor_5_a0_combout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_186_a21_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_186_a21.extended_lut = "off";
defparam fp_functions_0_aMux_186_a21.lut_mask = 64'h220A220A220A220A;
defparam fp_functions_0_aMux_186_a21.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai3365_a9(
	.dataa(!fp_functions_0_aMux_186_a11_combout),
	.datab(!fp_functions_0_aMux_186_a19_combout),
	.datac(!fp_functions_0_aMux_186_a13_combout),
	.datad(!fp_functions_0_aMux_186_a21_combout),
	.datae(!fp_functions_0_areduce_nor_4_acombout),
	.dataf(!fp_functions_0_arVStage_uid177_lzCountVal_uid85_fpAddTest_b_a0_a_a1_combout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai3365_a9_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai3365_a9.extended_lut = "off";
defparam fp_functions_0_ai3365_a9.lut_mask = 64'h0F0F00FF55553333;
defparam fp_functions_0_ai3365_a9.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_186_a22(
	.dataa(!fp_functions_0_aredist0_vStage_uid154_lzCountVal_uid85_fpAddTest_b_1_q_a7_a_aq),
	.datab(!fp_functions_0_aredist3_fracGRS_uid84_fpAddTest_q_1_q_a15_a_aq),
	.datac(!fp_functions_0_areduce_nor_3_acombout),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_186_a22_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_186_a22.extended_lut = "off";
defparam fp_functions_0_aMux_186_a22.lut_mask = 64'h5353535353535353;
defparam fp_functions_0_aMux_186_a22.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_186_a23(
	.dataa(!fp_functions_0_aredist1_vCount_uid152_lzCountVal_uid85_fpAddTest_q_1_q_a0_a_aq),
	.datab(!fp_functions_0_aMux_186_a18_combout),
	.datac(!fp_functions_0_aMux_186_a22_combout),
	.datad(!fp_functions_0_areduce_nor_5_a0_combout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_186_a23_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_186_a23.extended_lut = "off";
defparam fp_functions_0_aMux_186_a23.lut_mask = 64'h220A220A220A220A;
defparam fp_functions_0_aMux_186_a23.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai3365_a10(
	.dataa(!fp_functions_0_aMux_186_a13_combout),
	.datab(!fp_functions_0_aMux_186_a21_combout),
	.datac(!fp_functions_0_aMux_186_a15_combout),
	.datad(!fp_functions_0_aMux_186_a23_combout),
	.datae(!fp_functions_0_areduce_nor_4_acombout),
	.dataf(!fp_functions_0_arVStage_uid177_lzCountVal_uid85_fpAddTest_b_a0_a_a1_combout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai3365_a10_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai3365_a10.extended_lut = "off";
defparam fp_functions_0_ai3365_a10.lut_mask = 64'h0F0F00FF55553333;
defparam fp_functions_0_ai3365_a10.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_158_a0(
	.dataa(!fp_functions_0_aredist1_vCount_uid152_lzCountVal_uid85_fpAddTest_q_1_q_a0_a_aq),
	.datab(!fp_functions_0_aredist0_vStage_uid154_lzCountVal_uid85_fpAddTest_b_1_q_a0_a_aq),
	.datac(!fp_functions_0_aredist0_vStage_uid154_lzCountVal_uid85_fpAddTest_b_1_q_a8_a_aq),
	.datad(!fp_functions_0_aredist3_fracGRS_uid84_fpAddTest_q_1_q_a16_a_aq),
	.datae(!fp_functions_0_areduce_nor_3_acombout),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_158_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_158_a0.extended_lut = "off";
defparam fp_functions_0_aMux_158_a0.lut_mask = 64'h0A0A11BB0A0A11BB;
defparam fp_functions_0_aMux_158_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_186_a24(
	.dataa(!fp_functions_0_aredist1_vCount_uid152_lzCountVal_uid85_fpAddTest_q_1_q_a0_a_aq),
	.datab(!fp_functions_0_aMux_186_a20_combout),
	.datac(!fp_functions_0_aMux_158_a0_combout),
	.datad(!fp_functions_0_areduce_nor_5_a0_combout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_186_a24_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_186_a24.extended_lut = "off";
defparam fp_functions_0_aMux_186_a24.lut_mask = 64'h220F220F220F220F;
defparam fp_functions_0_aMux_186_a24.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai3365_a11(
	.dataa(!fp_functions_0_aMux_186_a15_combout),
	.datab(!fp_functions_0_aMux_186_a23_combout),
	.datac(!fp_functions_0_aMux_186_a17_combout),
	.datad(!fp_functions_0_aMux_186_a24_combout),
	.datae(!fp_functions_0_areduce_nor_4_acombout),
	.dataf(!fp_functions_0_arVStage_uid177_lzCountVal_uid85_fpAddTest_b_a0_a_a1_combout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai3365_a11_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai3365_a11.extended_lut = "off";
defparam fp_functions_0_ai3365_a11.lut_mask = 64'h0F0F00FF55553333;
defparam fp_functions_0_ai3365_a11.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_158_a1(
	.dataa(!fp_functions_0_aredist1_vCount_uid152_lzCountVal_uid85_fpAddTest_q_1_q_a0_a_aq),
	.datab(!fp_functions_0_aredist0_vStage_uid154_lzCountVal_uid85_fpAddTest_b_1_q_a1_a_aq),
	.datac(!fp_functions_0_aredist0_vStage_uid154_lzCountVal_uid85_fpAddTest_b_1_q_a9_a_aq),
	.datad(!fp_functions_0_aredist3_fracGRS_uid84_fpAddTest_q_1_q_a17_a_aq),
	.datae(!fp_functions_0_areduce_nor_3_acombout),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_158_a1_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_158_a1.extended_lut = "off";
defparam fp_functions_0_aMux_158_a1.lut_mask = 64'h0A0A11BB0A0A11BB;
defparam fp_functions_0_aMux_158_a1.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_186_a25(
	.dataa(!fp_functions_0_aredist1_vCount_uid152_lzCountVal_uid85_fpAddTest_q_1_q_a0_a_aq),
	.datab(!fp_functions_0_aMux_186_a22_combout),
	.datac(!fp_functions_0_aMux_158_a1_combout),
	.datad(!fp_functions_0_areduce_nor_5_a0_combout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_186_a25_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_186_a25.extended_lut = "off";
defparam fp_functions_0_aMux_186_a25.lut_mask = 64'h220F220F220F220F;
defparam fp_functions_0_aMux_186_a25.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai3365_a12(
	.dataa(!fp_functions_0_aMux_186_a17_combout),
	.datab(!fp_functions_0_aMux_186_a24_combout),
	.datac(!fp_functions_0_aMux_186_a19_combout),
	.datad(!fp_functions_0_aMux_186_a25_combout),
	.datae(!fp_functions_0_areduce_nor_4_acombout),
	.dataf(!fp_functions_0_arVStage_uid177_lzCountVal_uid85_fpAddTest_b_a0_a_a1_combout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai3365_a12_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai3365_a12.extended_lut = "off";
defparam fp_functions_0_ai3365_a12.lut_mask = 64'h0F0F00FF55553333;
defparam fp_functions_0_ai3365_a12.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_158_a2(
	.dataa(!fp_functions_0_aredist1_vCount_uid152_lzCountVal_uid85_fpAddTest_q_1_q_a0_a_aq),
	.datab(!fp_functions_0_aredist0_vStage_uid154_lzCountVal_uid85_fpAddTest_b_1_q_a2_a_aq),
	.datac(!fp_functions_0_aredist0_vStage_uid154_lzCountVal_uid85_fpAddTest_b_1_q_a10_a_aq),
	.datad(!fp_functions_0_aredist3_fracGRS_uid84_fpAddTest_q_1_q_a18_a_aq),
	.datae(!fp_functions_0_areduce_nor_3_acombout),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_158_a2_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_158_a2.extended_lut = "off";
defparam fp_functions_0_aMux_158_a2.lut_mask = 64'h0A0A11BB0A0A11BB;
defparam fp_functions_0_aMux_158_a2.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_186_a26(
	.dataa(!fp_functions_0_aMux_158_a0_combout),
	.datab(!fp_functions_0_aMux_158_a2_combout),
	.datac(!fp_functions_0_areduce_nor_5_a0_combout),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_186_a26_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_186_a26.extended_lut = "off";
defparam fp_functions_0_aMux_186_a26.lut_mask = 64'h5353535353535353;
defparam fp_functions_0_aMux_186_a26.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai3365_a13(
	.dataa(!fp_functions_0_aMux_186_a19_combout),
	.datab(!fp_functions_0_aMux_186_a25_combout),
	.datac(!fp_functions_0_aMux_186_a21_combout),
	.datad(!fp_functions_0_aMux_186_a26_combout),
	.datae(!fp_functions_0_areduce_nor_4_acombout),
	.dataf(!fp_functions_0_arVStage_uid177_lzCountVal_uid85_fpAddTest_b_a0_a_a1_combout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai3365_a13_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai3365_a13.extended_lut = "off";
defparam fp_functions_0_ai3365_a13.lut_mask = 64'h0F0F00FF55553333;
defparam fp_functions_0_ai3365_a13.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_158_a3(
	.dataa(!fp_functions_0_aredist1_vCount_uid152_lzCountVal_uid85_fpAddTest_q_1_q_a0_a_aq),
	.datab(!fp_functions_0_aredist0_vStage_uid154_lzCountVal_uid85_fpAddTest_b_1_q_a3_a_aq),
	.datac(!fp_functions_0_aredist3_fracGRS_uid84_fpAddTest_q_1_q_a11_a_aq),
	.datad(!fp_functions_0_aredist3_fracGRS_uid84_fpAddTest_q_1_q_a19_a_aq),
	.datae(!fp_functions_0_areduce_nor_3_acombout),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_158_a3_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_158_a3.extended_lut = "off";
defparam fp_functions_0_aMux_158_a3.lut_mask = 64'h0A0A11BB0A0A11BB;
defparam fp_functions_0_aMux_158_a3.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_186_a27(
	.dataa(!fp_functions_0_aMux_158_a1_combout),
	.datab(!fp_functions_0_aMux_158_a3_combout),
	.datac(!fp_functions_0_areduce_nor_5_a0_combout),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_186_a27_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_186_a27.extended_lut = "off";
defparam fp_functions_0_aMux_186_a27.lut_mask = 64'h5353535353535353;
defparam fp_functions_0_aMux_186_a27.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai3365_a14(
	.dataa(!fp_functions_0_aMux_186_a21_combout),
	.datab(!fp_functions_0_aMux_186_a26_combout),
	.datac(!fp_functions_0_aMux_186_a23_combout),
	.datad(!fp_functions_0_aMux_186_a27_combout),
	.datae(!fp_functions_0_areduce_nor_4_acombout),
	.dataf(!fp_functions_0_arVStage_uid177_lzCountVal_uid85_fpAddTest_b_a0_a_a1_combout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai3365_a14_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai3365_a14.extended_lut = "off";
defparam fp_functions_0_ai3365_a14.lut_mask = 64'h0F0F00FF55553333;
defparam fp_functions_0_ai3365_a14.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_158_a4(
	.dataa(!fp_functions_0_aredist1_vCount_uid152_lzCountVal_uid85_fpAddTest_q_1_q_a0_a_aq),
	.datab(!fp_functions_0_aredist0_vStage_uid154_lzCountVal_uid85_fpAddTest_b_1_q_a4_a_aq),
	.datac(!fp_functions_0_aredist3_fracGRS_uid84_fpAddTest_q_1_q_a12_a_aq),
	.datad(!fp_functions_0_aredist3_fracGRS_uid84_fpAddTest_q_1_q_a20_a_aq),
	.datae(!fp_functions_0_areduce_nor_3_acombout),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_158_a4_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_158_a4.extended_lut = "off";
defparam fp_functions_0_aMux_158_a4.lut_mask = 64'h0A0A11BB0A0A11BB;
defparam fp_functions_0_aMux_158_a4.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_186_a28(
	.dataa(!fp_functions_0_aMux_158_a2_combout),
	.datab(!fp_functions_0_aMux_158_a4_combout),
	.datac(!fp_functions_0_areduce_nor_5_a0_combout),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_186_a28_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_186_a28.extended_lut = "off";
defparam fp_functions_0_aMux_186_a28.lut_mask = 64'h5353535353535353;
defparam fp_functions_0_aMux_186_a28.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai3365_a15(
	.dataa(!fp_functions_0_aMux_186_a23_combout),
	.datab(!fp_functions_0_aMux_186_a27_combout),
	.datac(!fp_functions_0_aMux_186_a24_combout),
	.datad(!fp_functions_0_aMux_186_a28_combout),
	.datae(!fp_functions_0_areduce_nor_4_acombout),
	.dataf(!fp_functions_0_arVStage_uid177_lzCountVal_uid85_fpAddTest_b_a0_a_a1_combout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai3365_a15_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai3365_a15.extended_lut = "off";
defparam fp_functions_0_ai3365_a15.lut_mask = 64'h0F0F00FF55553333;
defparam fp_functions_0_ai3365_a15.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_158_a5(
	.dataa(!fp_functions_0_aredist1_vCount_uid152_lzCountVal_uid85_fpAddTest_q_1_q_a0_a_aq),
	.datab(!fp_functions_0_aredist0_vStage_uid154_lzCountVal_uid85_fpAddTest_b_1_q_a5_a_aq),
	.datac(!fp_functions_0_aredist3_fracGRS_uid84_fpAddTest_q_1_q_a13_a_aq),
	.datad(!fp_functions_0_aredist3_fracGRS_uid84_fpAddTest_q_1_q_a21_a_aq),
	.datae(!fp_functions_0_areduce_nor_3_acombout),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_158_a5_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_158_a5.extended_lut = "off";
defparam fp_functions_0_aMux_158_a5.lut_mask = 64'h0A0A11BB0A0A11BB;
defparam fp_functions_0_aMux_158_a5.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_186_a29(
	.dataa(!fp_functions_0_aMux_158_a3_combout),
	.datab(!fp_functions_0_aMux_158_a5_combout),
	.datac(!fp_functions_0_areduce_nor_5_a0_combout),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_186_a29_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_186_a29.extended_lut = "off";
defparam fp_functions_0_aMux_186_a29.lut_mask = 64'h5353535353535353;
defparam fp_functions_0_aMux_186_a29.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai3365_a16(
	.dataa(!fp_functions_0_aMux_186_a24_combout),
	.datab(!fp_functions_0_aMux_186_a28_combout),
	.datac(!fp_functions_0_aMux_186_a25_combout),
	.datad(!fp_functions_0_aMux_186_a29_combout),
	.datae(!fp_functions_0_areduce_nor_4_acombout),
	.dataf(!fp_functions_0_arVStage_uid177_lzCountVal_uid85_fpAddTest_b_a0_a_a1_combout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai3365_a16_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai3365_a16.extended_lut = "off";
defparam fp_functions_0_ai3365_a16.lut_mask = 64'h0F0F00FF55553333;
defparam fp_functions_0_ai3365_a16.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_158_a6(
	.dataa(!fp_functions_0_aredist1_vCount_uid152_lzCountVal_uid85_fpAddTest_q_1_q_a0_a_aq),
	.datab(!fp_functions_0_aredist0_vStage_uid154_lzCountVal_uid85_fpAddTest_b_1_q_a6_a_aq),
	.datac(!fp_functions_0_aredist3_fracGRS_uid84_fpAddTest_q_1_q_a14_a_aq),
	.datad(!fp_functions_0_aredist3_fracGRS_uid84_fpAddTest_q_1_q_a22_a_aq),
	.datae(!fp_functions_0_areduce_nor_3_acombout),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_158_a6_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_158_a6.extended_lut = "off";
defparam fp_functions_0_aMux_158_a6.lut_mask = 64'h0A0A11BB0A0A11BB;
defparam fp_functions_0_aMux_158_a6.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_186_a30(
	.dataa(!fp_functions_0_aMux_158_a4_combout),
	.datab(!fp_functions_0_aMux_158_a6_combout),
	.datac(!fp_functions_0_areduce_nor_5_a0_combout),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_186_a30_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_186_a30.extended_lut = "off";
defparam fp_functions_0_aMux_186_a30.lut_mask = 64'h5353535353535353;
defparam fp_functions_0_aMux_186_a30.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai3365_a17(
	.dataa(!fp_functions_0_aMux_186_a25_combout),
	.datab(!fp_functions_0_aMux_186_a29_combout),
	.datac(!fp_functions_0_aMux_186_a26_combout),
	.datad(!fp_functions_0_aMux_186_a30_combout),
	.datae(!fp_functions_0_areduce_nor_4_acombout),
	.dataf(!fp_functions_0_arVStage_uid177_lzCountVal_uid85_fpAddTest_b_a0_a_a1_combout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai3365_a17_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai3365_a17.extended_lut = "off";
defparam fp_functions_0_ai3365_a17.lut_mask = 64'h0F0F00FF55553333;
defparam fp_functions_0_ai3365_a17.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_158_a7(
	.dataa(!fp_functions_0_aredist1_vCount_uid152_lzCountVal_uid85_fpAddTest_q_1_q_a0_a_aq),
	.datab(!fp_functions_0_aredist0_vStage_uid154_lzCountVal_uid85_fpAddTest_b_1_q_a7_a_aq),
	.datac(!fp_functions_0_aredist3_fracGRS_uid84_fpAddTest_q_1_q_a15_a_aq),
	.datad(!fp_functions_0_aredist3_fracGRS_uid84_fpAddTest_q_1_q_a23_a_aq),
	.datae(!fp_functions_0_areduce_nor_3_acombout),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_158_a7_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_158_a7.extended_lut = "off";
defparam fp_functions_0_aMux_158_a7.lut_mask = 64'h0A0A11BB0A0A11BB;
defparam fp_functions_0_aMux_158_a7.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_186_a31(
	.dataa(!fp_functions_0_aMux_158_a1_combout),
	.datab(!fp_functions_0_aMux_158_a3_combout),
	.datac(!fp_functions_0_aMux_158_a5_combout),
	.datad(!fp_functions_0_aMux_158_a7_combout),
	.datae(!fp_functions_0_areduce_nor_5_a0_combout),
	.dataf(!fp_functions_0_areduce_nor_4_acombout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_186_a31_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_186_a31.extended_lut = "off";
defparam fp_functions_0_aMux_186_a31.lut_mask = 64'h555533330F0F00FF;
defparam fp_functions_0_aMux_186_a31.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai3337_a1(
	.dataa(!fp_functions_0_areduce_nor_4_acombout),
	.datab(!fp_functions_0_aMux_186_a31_combout),
	.datac(!fp_functions_0_arVStage_uid177_lzCountVal_uid85_fpAddTest_b_a0_a_a1_combout),
	.datad(!fp_functions_0_aMux_186_a26_combout),
	.datae(!fp_functions_0_aMux_186_a30_combout),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai3337_a1_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai3337_a1.extended_lut = "off";
defparam fp_functions_0_ai3337_a1.lut_mask = 64'h303A353F303A353F;
defparam fp_functions_0_ai3337_a1.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_158_a8(
	.dataa(!fp_functions_0_aredist3_fracGRS_uid84_fpAddTest_q_1_q_a16_a_aq),
	.datab(!fp_functions_0_aredist3_fracGRS_uid84_fpAddTest_q_1_q_a24_a_aq),
	.datac(!fp_functions_0_aredist0_vStage_uid154_lzCountVal_uid85_fpAddTest_b_1_q_a0_a_aq),
	.datad(!fp_functions_0_aredist0_vStage_uid154_lzCountVal_uid85_fpAddTest_b_1_q_a8_a_aq),
	.datae(!fp_functions_0_areduce_nor_3_acombout),
	.dataf(!fp_functions_0_aredist1_vCount_uid152_lzCountVal_uid85_fpAddTest_q_1_q_a0_a_aq),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_158_a8_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_158_a8.extended_lut = "off";
defparam fp_functions_0_aMux_158_a8.lut_mask = 64'h555533330F0F00FF;
defparam fp_functions_0_aMux_158_a8.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_186_a32(
	.dataa(!fp_functions_0_aMux_158_a2_combout),
	.datab(!fp_functions_0_aMux_158_a4_combout),
	.datac(!fp_functions_0_aMux_158_a6_combout),
	.datad(!fp_functions_0_aMux_158_a8_combout),
	.datae(!fp_functions_0_areduce_nor_5_a0_combout),
	.dataf(!fp_functions_0_areduce_nor_4_acombout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_186_a32_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_186_a32.extended_lut = "off";
defparam fp_functions_0_aMux_186_a32.lut_mask = 64'h555533330F0F00FF;
defparam fp_functions_0_aMux_186_a32.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai3365_a18(
	.dataa(!fp_functions_0_aMux_186_a31_combout),
	.datab(!fp_functions_0_aMux_186_a32_combout),
	.datac(!fp_functions_0_arVStage_uid177_lzCountVal_uid85_fpAddTest_b_a0_a_a1_combout),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai3365_a18_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai3365_a18.extended_lut = "off";
defparam fp_functions_0_ai3365_a18.lut_mask = 64'h3535353535353535;
defparam fp_functions_0_ai3365_a18.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_158_a9(
	.dataa(!fp_functions_0_aredist3_fracGRS_uid84_fpAddTest_q_1_q_a17_a_aq),
	.datab(!fp_functions_0_aredist3_fracGRS_uid84_fpAddTest_q_1_q_a25_a_aq),
	.datac(!fp_functions_0_aredist0_vStage_uid154_lzCountVal_uid85_fpAddTest_b_1_q_a1_a_aq),
	.datad(!fp_functions_0_aredist0_vStage_uid154_lzCountVal_uid85_fpAddTest_b_1_q_a9_a_aq),
	.datae(!fp_functions_0_areduce_nor_3_acombout),
	.dataf(!fp_functions_0_aredist1_vCount_uid152_lzCountVal_uid85_fpAddTest_q_1_q_a0_a_aq),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_158_a9_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_158_a9.extended_lut = "off";
defparam fp_functions_0_aMux_158_a9.lut_mask = 64'h555533330F0F00FF;
defparam fp_functions_0_aMux_158_a9.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_186_a33(
	.dataa(!fp_functions_0_aMux_158_a3_combout),
	.datab(!fp_functions_0_aMux_158_a5_combout),
	.datac(!fp_functions_0_aMux_158_a7_combout),
	.datad(!fp_functions_0_aMux_158_a9_combout),
	.datae(!fp_functions_0_areduce_nor_5_a0_combout),
	.dataf(!fp_functions_0_areduce_nor_4_acombout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_186_a33_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_186_a33.extended_lut = "off";
defparam fp_functions_0_aMux_186_a33.lut_mask = 64'h555533330F0F00FF;
defparam fp_functions_0_aMux_186_a33.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai3365_a19(
	.dataa(!fp_functions_0_aMux_186_a32_combout),
	.datab(!fp_functions_0_aMux_186_a33_combout),
	.datac(!fp_functions_0_arVStage_uid177_lzCountVal_uid85_fpAddTest_b_a0_a_a1_combout),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai3365_a19_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai3365_a19.extended_lut = "off";
defparam fp_functions_0_ai3365_a19.lut_mask = 64'h3535353535353535;
defparam fp_functions_0_ai3365_a19.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_158_a10(
	.dataa(!fp_functions_0_aredist3_fracGRS_uid84_fpAddTest_q_1_q_a18_a_aq),
	.datab(!fp_functions_0_aredist3_fracGRS_uid84_fpAddTest_q_1_q_a26_a_aq),
	.datac(!fp_functions_0_aredist0_vStage_uid154_lzCountVal_uid85_fpAddTest_b_1_q_a2_a_aq),
	.datad(!fp_functions_0_aredist0_vStage_uid154_lzCountVal_uid85_fpAddTest_b_1_q_a10_a_aq),
	.datae(!fp_functions_0_areduce_nor_3_acombout),
	.dataf(!fp_functions_0_aredist1_vCount_uid152_lzCountVal_uid85_fpAddTest_q_1_q_a0_a_aq),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_158_a10_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_158_a10.extended_lut = "off";
defparam fp_functions_0_aMux_158_a10.lut_mask = 64'h555533330F0F00FF;
defparam fp_functions_0_aMux_158_a10.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_186_a34(
	.dataa(!fp_functions_0_aMux_158_a4_combout),
	.datab(!fp_functions_0_aMux_158_a6_combout),
	.datac(!fp_functions_0_aMux_158_a8_combout),
	.datad(!fp_functions_0_aMux_158_a10_combout),
	.datae(!fp_functions_0_areduce_nor_5_a0_combout),
	.dataf(!fp_functions_0_areduce_nor_4_acombout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_186_a34_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_186_a34.extended_lut = "off";
defparam fp_functions_0_aMux_186_a34.lut_mask = 64'h555533330F0F00FF;
defparam fp_functions_0_aMux_186_a34.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai3337_a2(
	.dataa(!fp_functions_0_aMux_186_a33_combout),
	.datab(!fp_functions_0_aMux_186_a34_combout),
	.datac(!fp_functions_0_arVStage_uid177_lzCountVal_uid85_fpAddTest_b_a0_a_a1_combout),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai3337_a2_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai3337_a2.extended_lut = "off";
defparam fp_functions_0_ai3337_a2.lut_mask = 64'h3535353535353535;
defparam fp_functions_0_ai3337_a2.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_astickyBits_uid69_fpAddTest_merged_bit_select_b_a0_a_a0(
	.dataa(!fp_functions_0_ashiftedOut_uid63_fpAddTest_o_a10_a_aq),
	.datab(!fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a42_a_aq),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_astickyBits_uid69_fpAddTest_merged_bit_select_b_a0_a_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_astickyBits_uid69_fpAddTest_merged_bit_select_b_a0_a_a0.extended_lut = "off";
defparam fp_functions_0_astickyBits_uid69_fpAddTest_merged_bit_select_b_a0_a_a0.lut_mask = 64'h2222222222222222;
defparam fp_functions_0_astickyBits_uid69_fpAddTest_merged_bit_select_b_a0_a_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_astickyBits_uid69_fpAddTest_merged_bit_select_b_a0_a_a1(
	.dataa(!fp_functions_0_ashiftedOut_uid63_fpAddTest_o_a10_a_aq),
	.datab(!fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a38_a_aq),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_astickyBits_uid69_fpAddTest_merged_bit_select_b_a0_a_a1_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_astickyBits_uid69_fpAddTest_merged_bit_select_b_a0_a_a1.extended_lut = "off";
defparam fp_functions_0_astickyBits_uid69_fpAddTest_merged_bit_select_b_a0_a_a1.lut_mask = 64'h2222222222222222;
defparam fp_functions_0_astickyBits_uid69_fpAddTest_merged_bit_select_b_a0_a_a1.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_astickyBits_uid69_fpAddTest_merged_bit_select_b_a0_a_a2(
	.dataa(!fp_functions_0_ashiftedOut_uid63_fpAddTest_o_a10_a_aq),
	.datab(!fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a34_a_aq),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_astickyBits_uid69_fpAddTest_merged_bit_select_b_a0_a_a2_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_astickyBits_uid69_fpAddTest_merged_bit_select_b_a0_a_a2.extended_lut = "off";
defparam fp_functions_0_astickyBits_uid69_fpAddTest_merged_bit_select_b_a0_a_a2.lut_mask = 64'h2222222222222222;
defparam fp_functions_0_astickyBits_uid69_fpAddTest_merged_bit_select_b_a0_a_a2.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_astickyBits_uid69_fpAddTest_merged_bit_select_b_a0_a_a3(
	.dataa(!fp_functions_0_ashiftedOut_uid63_fpAddTest_o_a10_a_aq),
	.datab(!fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a35_a_aq),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_astickyBits_uid69_fpAddTest_merged_bit_select_b_a0_a_a3_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_astickyBits_uid69_fpAddTest_merged_bit_select_b_a0_a_a3.extended_lut = "off";
defparam fp_functions_0_astickyBits_uid69_fpAddTest_merged_bit_select_b_a0_a_a3.lut_mask = 64'h2222222222222222;
defparam fp_functions_0_astickyBits_uid69_fpAddTest_merged_bit_select_b_a0_a_a3.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_astickyBits_uid69_fpAddTest_merged_bit_select_b_a0_a_a4(
	.dataa(!fp_functions_0_ashiftedOut_uid63_fpAddTest_o_a10_a_aq),
	.datab(!fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a36_a_aq),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_astickyBits_uid69_fpAddTest_merged_bit_select_b_a0_a_a4_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_astickyBits_uid69_fpAddTest_merged_bit_select_b_a0_a_a4.extended_lut = "off";
defparam fp_functions_0_astickyBits_uid69_fpAddTest_merged_bit_select_b_a0_a_a4.lut_mask = 64'h2222222222222222;
defparam fp_functions_0_astickyBits_uid69_fpAddTest_merged_bit_select_b_a0_a_a4.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_astickyBits_uid69_fpAddTest_merged_bit_select_b_a0_a_a5(
	.dataa(!fp_functions_0_ashiftedOut_uid63_fpAddTest_o_a10_a_aq),
	.datab(!fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a37_a_aq),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_astickyBits_uid69_fpAddTest_merged_bit_select_b_a0_a_a5_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_astickyBits_uid69_fpAddTest_merged_bit_select_b_a0_a_a5.extended_lut = "off";
defparam fp_functions_0_astickyBits_uid69_fpAddTest_merged_bit_select_b_a0_a_a5.lut_mask = 64'h2222222222222222;
defparam fp_functions_0_astickyBits_uid69_fpAddTest_merged_bit_select_b_a0_a_a5.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_astickyBits_uid69_fpAddTest_merged_bit_select_b_a0_a_a6(
	.dataa(!fp_functions_0_ashiftedOut_uid63_fpAddTest_o_a10_a_aq),
	.datab(!fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a39_a_aq),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_astickyBits_uid69_fpAddTest_merged_bit_select_b_a0_a_a6_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_astickyBits_uid69_fpAddTest_merged_bit_select_b_a0_a_a6.extended_lut = "off";
defparam fp_functions_0_astickyBits_uid69_fpAddTest_merged_bit_select_b_a0_a_a6.lut_mask = 64'h2222222222222222;
defparam fp_functions_0_astickyBits_uid69_fpAddTest_merged_bit_select_b_a0_a_a6.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_astickyBits_uid69_fpAddTest_merged_bit_select_b_a0_a_a7(
	.dataa(!fp_functions_0_ashiftedOut_uid63_fpAddTest_o_a10_a_aq),
	.datab(!fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a40_a_aq),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_astickyBits_uid69_fpAddTest_merged_bit_select_b_a0_a_a7_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_astickyBits_uid69_fpAddTest_merged_bit_select_b_a0_a_a7.extended_lut = "off";
defparam fp_functions_0_astickyBits_uid69_fpAddTest_merged_bit_select_b_a0_a_a7.lut_mask = 64'h2222222222222222;
defparam fp_functions_0_astickyBits_uid69_fpAddTest_merged_bit_select_b_a0_a_a7.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_astickyBits_uid69_fpAddTest_merged_bit_select_b_a0_a_a8(
	.dataa(!fp_functions_0_ashiftedOut_uid63_fpAddTest_o_a10_a_aq),
	.datab(!fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a41_a_aq),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_astickyBits_uid69_fpAddTest_merged_bit_select_b_a0_a_a8_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_astickyBits_uid69_fpAddTest_merged_bit_select_b_a0_a_a8.extended_lut = "off";
defparam fp_functions_0_astickyBits_uid69_fpAddTest_merged_bit_select_b_a0_a_a8.lut_mask = 64'h2222222222222222;
defparam fp_functions_0_astickyBits_uid69_fpAddTest_merged_bit_select_b_a0_a_a8.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_astickyBits_uid69_fpAddTest_merged_bit_select_b_a0_a_a9(
	.dataa(!fp_functions_0_ashiftedOut_uid63_fpAddTest_o_a10_a_aq),
	.datab(!fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a47_a_aq),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_astickyBits_uid69_fpAddTest_merged_bit_select_b_a0_a_a9_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_astickyBits_uid69_fpAddTest_merged_bit_select_b_a0_a_a9.extended_lut = "off";
defparam fp_functions_0_astickyBits_uid69_fpAddTest_merged_bit_select_b_a0_a_a9.lut_mask = 64'h2222222222222222;
defparam fp_functions_0_astickyBits_uid69_fpAddTest_merged_bit_select_b_a0_a_a9.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_astickyBits_uid69_fpAddTest_merged_bit_select_b_a0_a_a10(
	.dataa(!fp_functions_0_ashiftedOut_uid63_fpAddTest_o_a10_a_aq),
	.datab(!fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a43_a_aq),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_astickyBits_uid69_fpAddTest_merged_bit_select_b_a0_a_a10_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_astickyBits_uid69_fpAddTest_merged_bit_select_b_a0_a_a10.extended_lut = "off";
defparam fp_functions_0_astickyBits_uid69_fpAddTest_merged_bit_select_b_a0_a_a10.lut_mask = 64'h2222222222222222;
defparam fp_functions_0_astickyBits_uid69_fpAddTest_merged_bit_select_b_a0_a_a10.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_astickyBits_uid69_fpAddTest_merged_bit_select_b_a0_a_a11(
	.dataa(!fp_functions_0_ashiftedOut_uid63_fpAddTest_o_a10_a_aq),
	.datab(!fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a44_a_aq),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_astickyBits_uid69_fpAddTest_merged_bit_select_b_a0_a_a11_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_astickyBits_uid69_fpAddTest_merged_bit_select_b_a0_a_a11.extended_lut = "off";
defparam fp_functions_0_astickyBits_uid69_fpAddTest_merged_bit_select_b_a0_a_a11.lut_mask = 64'h2222222222222222;
defparam fp_functions_0_astickyBits_uid69_fpAddTest_merged_bit_select_b_a0_a_a11.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_astickyBits_uid69_fpAddTest_merged_bit_select_b_a0_a_a12(
	.dataa(!fp_functions_0_ashiftedOut_uid63_fpAddTest_o_a10_a_aq),
	.datab(!fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a45_a_aq),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_astickyBits_uid69_fpAddTest_merged_bit_select_b_a0_a_a12_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_astickyBits_uid69_fpAddTest_merged_bit_select_b_a0_a_a12.extended_lut = "off";
defparam fp_functions_0_astickyBits_uid69_fpAddTest_merged_bit_select_b_a0_a_a12.lut_mask = 64'h2222222222222222;
defparam fp_functions_0_astickyBits_uid69_fpAddTest_merged_bit_select_b_a0_a_a12.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_astickyBits_uid69_fpAddTest_merged_bit_select_b_a0_a_a13(
	.dataa(!fp_functions_0_ashiftedOut_uid63_fpAddTest_o_a10_a_aq),
	.datab(!fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a46_a_aq),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_astickyBits_uid69_fpAddTest_merged_bit_select_b_a0_a_a13_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_astickyBits_uid69_fpAddTest_merged_bit_select_b_a0_a_a13.extended_lut = "off";
defparam fp_functions_0_astickyBits_uid69_fpAddTest_merged_bit_select_b_a0_a_a13.lut_mask = 64'h2222222222222222;
defparam fp_functions_0_astickyBits_uid69_fpAddTest_merged_bit_select_b_a0_a_a13.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_astickyBits_uid69_fpAddTest_merged_bit_select_b_a0_a_a14(
	.dataa(!fp_functions_0_ashiftedOut_uid63_fpAddTest_o_a10_a_aq),
	.datab(!fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a29_a_aq),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_astickyBits_uid69_fpAddTest_merged_bit_select_b_a0_a_a14_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_astickyBits_uid69_fpAddTest_merged_bit_select_b_a0_a_a14.extended_lut = "off";
defparam fp_functions_0_astickyBits_uid69_fpAddTest_merged_bit_select_b_a0_a_a14.lut_mask = 64'h2222222222222222;
defparam fp_functions_0_astickyBits_uid69_fpAddTest_merged_bit_select_b_a0_a_a14.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_astickyBits_uid69_fpAddTest_merged_bit_select_b_a0_a_a15(
	.dataa(!fp_functions_0_ashiftedOut_uid63_fpAddTest_o_a10_a_aq),
	.datab(!fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a28_a_aq),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_astickyBits_uid69_fpAddTest_merged_bit_select_b_a0_a_a15_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_astickyBits_uid69_fpAddTest_merged_bit_select_b_a0_a_a15.extended_lut = "off";
defparam fp_functions_0_astickyBits_uid69_fpAddTest_merged_bit_select_b_a0_a_a15.lut_mask = 64'h2222222222222222;
defparam fp_functions_0_astickyBits_uid69_fpAddTest_merged_bit_select_b_a0_a_a15.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_astickyBits_uid69_fpAddTest_merged_bit_select_b_a0_a_a16(
	.dataa(!fp_functions_0_ashiftedOut_uid63_fpAddTest_o_a10_a_aq),
	.datab(!fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a26_a_aq),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_astickyBits_uid69_fpAddTest_merged_bit_select_b_a0_a_a16_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_astickyBits_uid69_fpAddTest_merged_bit_select_b_a0_a_a16.extended_lut = "off";
defparam fp_functions_0_astickyBits_uid69_fpAddTest_merged_bit_select_b_a0_a_a16.lut_mask = 64'h2222222222222222;
defparam fp_functions_0_astickyBits_uid69_fpAddTest_merged_bit_select_b_a0_a_a16.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_astickyBits_uid69_fpAddTest_merged_bit_select_b_a0_a_a17(
	.dataa(!fp_functions_0_ashiftedOut_uid63_fpAddTest_o_a10_a_aq),
	.datab(!fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a27_a_aq),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_astickyBits_uid69_fpAddTest_merged_bit_select_b_a0_a_a17_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_astickyBits_uid69_fpAddTest_merged_bit_select_b_a0_a_a17.extended_lut = "off";
defparam fp_functions_0_astickyBits_uid69_fpAddTest_merged_bit_select_b_a0_a_a17.lut_mask = 64'h2222222222222222;
defparam fp_functions_0_astickyBits_uid69_fpAddTest_merged_bit_select_b_a0_a_a17.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_astickyBits_uid69_fpAddTest_merged_bit_select_b_a0_a_a18(
	.dataa(!fp_functions_0_ashiftedOut_uid63_fpAddTest_o_a10_a_aq),
	.datab(!fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a33_a_aq),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_astickyBits_uid69_fpAddTest_merged_bit_select_b_a0_a_a18_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_astickyBits_uid69_fpAddTest_merged_bit_select_b_a0_a_a18.extended_lut = "off";
defparam fp_functions_0_astickyBits_uid69_fpAddTest_merged_bit_select_b_a0_a_a18.lut_mask = 64'h2222222222222222;
defparam fp_functions_0_astickyBits_uid69_fpAddTest_merged_bit_select_b_a0_a_a18.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_astickyBits_uid69_fpAddTest_merged_bit_select_b_a0_a_a19(
	.dataa(!fp_functions_0_ashiftedOut_uid63_fpAddTest_o_a10_a_aq),
	.datab(!fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a32_a_aq),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_astickyBits_uid69_fpAddTest_merged_bit_select_b_a0_a_a19_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_astickyBits_uid69_fpAddTest_merged_bit_select_b_a0_a_a19.extended_lut = "off";
defparam fp_functions_0_astickyBits_uid69_fpAddTest_merged_bit_select_b_a0_a_a19.lut_mask = 64'h2222222222222222;
defparam fp_functions_0_astickyBits_uid69_fpAddTest_merged_bit_select_b_a0_a_a19.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_astickyBits_uid69_fpAddTest_merged_bit_select_b_a0_a_a20(
	.dataa(!fp_functions_0_ashiftedOut_uid63_fpAddTest_o_a10_a_aq),
	.datab(!fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a25_a_aq),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_astickyBits_uid69_fpAddTest_merged_bit_select_b_a0_a_a20_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_astickyBits_uid69_fpAddTest_merged_bit_select_b_a0_a_a20.extended_lut = "off";
defparam fp_functions_0_astickyBits_uid69_fpAddTest_merged_bit_select_b_a0_a_a20.lut_mask = 64'h2222222222222222;
defparam fp_functions_0_astickyBits_uid69_fpAddTest_merged_bit_select_b_a0_a_a20.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_astickyBits_uid69_fpAddTest_merged_bit_select_b_a0_a_a21(
	.dataa(!fp_functions_0_ashiftedOut_uid63_fpAddTest_o_a10_a_aq),
	.datab(!fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a30_a_aq),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_astickyBits_uid69_fpAddTest_merged_bit_select_b_a0_a_a21_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_astickyBits_uid69_fpAddTest_merged_bit_select_b_a0_a_a21.extended_lut = "off";
defparam fp_functions_0_astickyBits_uid69_fpAddTest_merged_bit_select_b_a0_a_a21.lut_mask = 64'h2222222222222222;
defparam fp_functions_0_astickyBits_uid69_fpAddTest_merged_bit_select_b_a0_a_a21.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_astickyBits_uid69_fpAddTest_merged_bit_select_b_a0_a_a22(
	.dataa(!fp_functions_0_ashiftedOut_uid63_fpAddTest_o_a10_a_aq),
	.datab(!fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a31_a_aq),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_astickyBits_uid69_fpAddTest_merged_bit_select_b_a0_a_a22_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_astickyBits_uid69_fpAddTest_merged_bit_select_b_a0_a_a22.extended_lut = "off";
defparam fp_functions_0_astickyBits_uid69_fpAddTest_merged_bit_select_b_a0_a_a22.lut_mask = 64'h2222222222222222;
defparam fp_functions_0_astickyBits_uid69_fpAddTest_merged_bit_select_b_a0_a_a22.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_astickyBits_uid69_fpAddTest_merged_bit_select_b_a0_a_a23(
	.dataa(!fp_functions_0_ashiftedOut_uid63_fpAddTest_o_a10_a_aq),
	.datab(!fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a23_a_aq),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_astickyBits_uid69_fpAddTest_merged_bit_select_b_a0_a_a23_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_astickyBits_uid69_fpAddTest_merged_bit_select_b_a0_a_a23.extended_lut = "off";
defparam fp_functions_0_astickyBits_uid69_fpAddTest_merged_bit_select_b_a0_a_a23.lut_mask = 64'h2222222222222222;
defparam fp_functions_0_astickyBits_uid69_fpAddTest_merged_bit_select_b_a0_a_a23.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_afrac_bSig_uid36_fpAddTest_b_a13_a_a0(
	.dataa(!b[13]),
	.datab(!a[13]),
	.datac(!fp_functions_0_aadd_0_a1_sumout),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_afrac_bSig_uid36_fpAddTest_b_a13_a_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_afrac_bSig_uid36_fpAddTest_b_a13_a_a0.extended_lut = "off";
defparam fp_functions_0_afrac_bSig_uid36_fpAddTest_b_a13_a_a0.lut_mask = 64'h5353535353535353;
defparam fp_functions_0_afrac_bSig_uid36_fpAddTest_b_a13_a_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_afrac_bSig_uid36_fpAddTest_b_a14_a_a1(
	.dataa(!b[14]),
	.datab(!a[14]),
	.datac(!fp_functions_0_aadd_0_a1_sumout),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_afrac_bSig_uid36_fpAddTest_b_a14_a_a1_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_afrac_bSig_uid36_fpAddTest_b_a14_a_a1.extended_lut = "off";
defparam fp_functions_0_afrac_bSig_uid36_fpAddTest_b_a14_a_a1.lut_mask = 64'h5353535353535353;
defparam fp_functions_0_afrac_bSig_uid36_fpAddTest_b_a14_a_a1.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_areduce_nor_0_a0(
	.dataa(!b[30]),
	.datab(!a[30]),
	.datac(!b[29]),
	.datad(!a[29]),
	.datae(!fp_functions_0_aadd_0_a1_sumout),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_areduce_nor_0_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_areduce_nor_0_a0.extended_lut = "off";
defparam fp_functions_0_areduce_nor_0_a0.lut_mask = 64'hA0A0CC00A0A0CC00;
defparam fp_functions_0_areduce_nor_0_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_areduce_nor_0_a1(
	.dataa(!b[28]),
	.datab(!a[28]),
	.datac(!b[27]),
	.datad(!a[27]),
	.datae(!fp_functions_0_aadd_0_a1_sumout),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_areduce_nor_0_a1_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_areduce_nor_0_a1.extended_lut = "off";
defparam fp_functions_0_areduce_nor_0_a1.lut_mask = 64'hA0A0CC00A0A0CC00;
defparam fp_functions_0_areduce_nor_0_a1.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_areduce_nor_0_a2(
	.dataa(!b[24]),
	.datab(!a[24]),
	.datac(!b[23]),
	.datad(!a[23]),
	.datae(!fp_functions_0_aadd_0_a1_sumout),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_areduce_nor_0_a2_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_areduce_nor_0_a2.extended_lut = "off";
defparam fp_functions_0_areduce_nor_0_a2.lut_mask = 64'hA0A0CC00A0A0CC00;
defparam fp_functions_0_areduce_nor_0_a2.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_areduce_nor_0_a3(
	.dataa(!b[26]),
	.datab(!a[26]),
	.datac(!b[25]),
	.datad(!a[25]),
	.datae(!fp_functions_0_aadd_0_a1_sumout),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_areduce_nor_0_a3_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_areduce_nor_0_a3.extended_lut = "off";
defparam fp_functions_0_areduce_nor_0_a3.lut_mask = 64'hA0A0CC00A0A0CC00;
defparam fp_functions_0_areduce_nor_0_a3.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_areduce_nor_0(
	.dataa(!fp_functions_0_areduce_nor_0_a0_combout),
	.datab(!fp_functions_0_areduce_nor_0_a1_combout),
	.datac(!fp_functions_0_areduce_nor_0_a2_combout),
	.datad(!fp_functions_0_areduce_nor_0_a3_combout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_areduce_nor_0_acombout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_areduce_nor_0.extended_lut = "off";
defparam fp_functions_0_areduce_nor_0.lut_mask = 64'hFFFEFFFEFFFEFFFE;
defparam fp_functions_0_areduce_nor_0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_2_a0(
	.dataa(!fp_functions_0_aadd_1_a11_sumout),
	.datab(!fp_functions_0_afrac_bSig_uid36_fpAddTest_b_a13_a_a0_combout),
	.datac(!fp_functions_0_afrac_bSig_uid36_fpAddTest_b_a14_a_a1_combout),
	.datad(!fp_functions_0_areduce_nor_0_acombout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_2_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_2_a0.extended_lut = "off";
defparam fp_functions_0_aMux_2_a0.lut_mask = 64'h0027002700270027;
defparam fp_functions_0_aMux_2_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_afrac_bSig_uid36_fpAddTest_b_a15_a_a2(
	.dataa(!b[15]),
	.datab(!a[15]),
	.datac(!fp_functions_0_aadd_0_a1_sumout),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_afrac_bSig_uid36_fpAddTest_b_a15_a_a2_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_afrac_bSig_uid36_fpAddTest_b_a15_a_a2.extended_lut = "off";
defparam fp_functions_0_afrac_bSig_uid36_fpAddTest_b_a15_a_a2.lut_mask = 64'h5353535353535353;
defparam fp_functions_0_afrac_bSig_uid36_fpAddTest_b_a15_a_a2.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_afrac_bSig_uid36_fpAddTest_b_a16_a_a3(
	.dataa(!b[16]),
	.datab(!a[16]),
	.datac(!fp_functions_0_aadd_0_a1_sumout),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_afrac_bSig_uid36_fpAddTest_b_a16_a_a3_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_afrac_bSig_uid36_fpAddTest_b_a16_a_a3.extended_lut = "off";
defparam fp_functions_0_afrac_bSig_uid36_fpAddTest_b_a16_a_a3.lut_mask = 64'h5353535353535353;
defparam fp_functions_0_afrac_bSig_uid36_fpAddTest_b_a16_a_a3.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_2_a1(
	.dataa(!fp_functions_0_aadd_1_a11_sumout),
	.datab(!fp_functions_0_afrac_bSig_uid36_fpAddTest_b_a15_a_a2_combout),
	.datac(!fp_functions_0_afrac_bSig_uid36_fpAddTest_b_a16_a_a3_combout),
	.datad(!fp_functions_0_areduce_nor_0_acombout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_2_a1_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_2_a1.extended_lut = "off";
defparam fp_functions_0_aMux_2_a1.lut_mask = 64'h0027002700270027;
defparam fp_functions_0_aMux_2_a1.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_afrac_bSig_uid36_fpAddTest_b_a17_a_a4(
	.dataa(!b[17]),
	.datab(!a[17]),
	.datac(!fp_functions_0_aadd_0_a1_sumout),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_afrac_bSig_uid36_fpAddTest_b_a17_a_a4_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_afrac_bSig_uid36_fpAddTest_b_a17_a_a4.extended_lut = "off";
defparam fp_functions_0_afrac_bSig_uid36_fpAddTest_b_a17_a_a4.lut_mask = 64'h5353535353535353;
defparam fp_functions_0_afrac_bSig_uid36_fpAddTest_b_a17_a_a4.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_afrac_bSig_uid36_fpAddTest_b_a18_a_a5(
	.dataa(!b[18]),
	.datab(!a[18]),
	.datac(!fp_functions_0_aadd_0_a1_sumout),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_afrac_bSig_uid36_fpAddTest_b_a18_a_a5_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_afrac_bSig_uid36_fpAddTest_b_a18_a_a5.extended_lut = "off";
defparam fp_functions_0_afrac_bSig_uid36_fpAddTest_b_a18_a_a5.lut_mask = 64'h5353535353535353;
defparam fp_functions_0_afrac_bSig_uid36_fpAddTest_b_a18_a_a5.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_2_a2(
	.dataa(!fp_functions_0_aadd_1_a11_sumout),
	.datab(!fp_functions_0_afrac_bSig_uid36_fpAddTest_b_a17_a_a4_combout),
	.datac(!fp_functions_0_afrac_bSig_uid36_fpAddTest_b_a18_a_a5_combout),
	.datad(!fp_functions_0_areduce_nor_0_acombout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_2_a2_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_2_a2.extended_lut = "off";
defparam fp_functions_0_aMux_2_a2.lut_mask = 64'h0027002700270027;
defparam fp_functions_0_aMux_2_a2.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_afrac_bSig_uid36_fpAddTest_b_a19_a_a6(
	.dataa(!b[19]),
	.datab(!a[19]),
	.datac(!fp_functions_0_aadd_0_a1_sumout),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_afrac_bSig_uid36_fpAddTest_b_a19_a_a6_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_afrac_bSig_uid36_fpAddTest_b_a19_a_a6.extended_lut = "off";
defparam fp_functions_0_afrac_bSig_uid36_fpAddTest_b_a19_a_a6.lut_mask = 64'h5353535353535353;
defparam fp_functions_0_afrac_bSig_uid36_fpAddTest_b_a19_a_a6.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_afrac_bSig_uid36_fpAddTest_b_a20_a_a7(
	.dataa(!b[20]),
	.datab(!a[20]),
	.datac(!fp_functions_0_aadd_0_a1_sumout),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_afrac_bSig_uid36_fpAddTest_b_a20_a_a7_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_afrac_bSig_uid36_fpAddTest_b_a20_a_a7.extended_lut = "off";
defparam fp_functions_0_afrac_bSig_uid36_fpAddTest_b_a20_a_a7.lut_mask = 64'h5353535353535353;
defparam fp_functions_0_afrac_bSig_uid36_fpAddTest_b_a20_a_a7.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_2_a3(
	.dataa(!fp_functions_0_aadd_1_a11_sumout),
	.datab(!fp_functions_0_afrac_bSig_uid36_fpAddTest_b_a19_a_a6_combout),
	.datac(!fp_functions_0_afrac_bSig_uid36_fpAddTest_b_a20_a_a7_combout),
	.datad(!fp_functions_0_areduce_nor_0_acombout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_2_a3_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_2_a3.extended_lut = "off";
defparam fp_functions_0_aMux_2_a3.lut_mask = 64'h0027002700270027;
defparam fp_functions_0_aMux_2_a3.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_59_a0(
	.dataa(!fp_functions_0_aMux_2_a0_combout),
	.datab(!fp_functions_0_aMux_2_a1_combout),
	.datac(!fp_functions_0_aMux_2_a2_combout),
	.datad(!fp_functions_0_aMux_2_a3_combout),
	.datae(!fp_functions_0_aadd_1_a16_sumout),
	.dataf(!fp_functions_0_aadd_1_a21_sumout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_59_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_59_a0.extended_lut = "off";
defparam fp_functions_0_aMux_59_a0.lut_mask = 64'h555533330F0F00FF;
defparam fp_functions_0_aMux_59_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_afrac_bSig_uid36_fpAddTest_b_a5_a_a8(
	.dataa(!b[5]),
	.datab(!a[5]),
	.datac(!fp_functions_0_aadd_0_a1_sumout),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_afrac_bSig_uid36_fpAddTest_b_a5_a_a8_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_afrac_bSig_uid36_fpAddTest_b_a5_a_a8.extended_lut = "off";
defparam fp_functions_0_afrac_bSig_uid36_fpAddTest_b_a5_a_a8.lut_mask = 64'h5353535353535353;
defparam fp_functions_0_afrac_bSig_uid36_fpAddTest_b_a5_a_a8.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_afrac_bSig_uid36_fpAddTest_b_a6_a_a9(
	.dataa(!b[6]),
	.datab(!a[6]),
	.datac(!fp_functions_0_aadd_0_a1_sumout),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_afrac_bSig_uid36_fpAddTest_b_a6_a_a9_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_afrac_bSig_uid36_fpAddTest_b_a6_a_a9.extended_lut = "off";
defparam fp_functions_0_afrac_bSig_uid36_fpAddTest_b_a6_a_a9.lut_mask = 64'h5353535353535353;
defparam fp_functions_0_afrac_bSig_uid36_fpAddTest_b_a6_a_a9.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_2_a4(
	.dataa(!fp_functions_0_aadd_1_a11_sumout),
	.datab(!fp_functions_0_afrac_bSig_uid36_fpAddTest_b_a5_a_a8_combout),
	.datac(!fp_functions_0_afrac_bSig_uid36_fpAddTest_b_a6_a_a9_combout),
	.datad(!fp_functions_0_areduce_nor_0_acombout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_2_a4_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_2_a4.extended_lut = "off";
defparam fp_functions_0_aMux_2_a4.lut_mask = 64'h0027002700270027;
defparam fp_functions_0_aMux_2_a4.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_afrac_bSig_uid36_fpAddTest_b_a7_a_a10(
	.dataa(!b[7]),
	.datab(!a[7]),
	.datac(!fp_functions_0_aadd_0_a1_sumout),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_afrac_bSig_uid36_fpAddTest_b_a7_a_a10_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_afrac_bSig_uid36_fpAddTest_b_a7_a_a10.extended_lut = "off";
defparam fp_functions_0_afrac_bSig_uid36_fpAddTest_b_a7_a_a10.lut_mask = 64'h5353535353535353;
defparam fp_functions_0_afrac_bSig_uid36_fpAddTest_b_a7_a_a10.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_afrac_bSig_uid36_fpAddTest_b_a8_a_a11(
	.dataa(!b[8]),
	.datab(!a[8]),
	.datac(!fp_functions_0_aadd_0_a1_sumout),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_afrac_bSig_uid36_fpAddTest_b_a8_a_a11_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_afrac_bSig_uid36_fpAddTest_b_a8_a_a11.extended_lut = "off";
defparam fp_functions_0_afrac_bSig_uid36_fpAddTest_b_a8_a_a11.lut_mask = 64'h5353535353535353;
defparam fp_functions_0_afrac_bSig_uid36_fpAddTest_b_a8_a_a11.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_2_a5(
	.dataa(!fp_functions_0_aadd_1_a11_sumout),
	.datab(!fp_functions_0_afrac_bSig_uid36_fpAddTest_b_a7_a_a10_combout),
	.datac(!fp_functions_0_afrac_bSig_uid36_fpAddTest_b_a8_a_a11_combout),
	.datad(!fp_functions_0_areduce_nor_0_acombout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_2_a5_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_2_a5.extended_lut = "off";
defparam fp_functions_0_aMux_2_a5.lut_mask = 64'h0027002700270027;
defparam fp_functions_0_aMux_2_a5.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_afrac_bSig_uid36_fpAddTest_b_a9_a_a12(
	.dataa(!b[9]),
	.datab(!a[9]),
	.datac(!fp_functions_0_aadd_0_a1_sumout),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_afrac_bSig_uid36_fpAddTest_b_a9_a_a12_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_afrac_bSig_uid36_fpAddTest_b_a9_a_a12.extended_lut = "off";
defparam fp_functions_0_afrac_bSig_uid36_fpAddTest_b_a9_a_a12.lut_mask = 64'h5353535353535353;
defparam fp_functions_0_afrac_bSig_uid36_fpAddTest_b_a9_a_a12.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_afrac_bSig_uid36_fpAddTest_b_a10_a_a13(
	.dataa(!b[10]),
	.datab(!a[10]),
	.datac(!fp_functions_0_aadd_0_a1_sumout),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_afrac_bSig_uid36_fpAddTest_b_a10_a_a13_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_afrac_bSig_uid36_fpAddTest_b_a10_a_a13.extended_lut = "off";
defparam fp_functions_0_afrac_bSig_uid36_fpAddTest_b_a10_a_a13.lut_mask = 64'h5353535353535353;
defparam fp_functions_0_afrac_bSig_uid36_fpAddTest_b_a10_a_a13.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_2_a6(
	.dataa(!fp_functions_0_aadd_1_a11_sumout),
	.datab(!fp_functions_0_afrac_bSig_uid36_fpAddTest_b_a9_a_a12_combout),
	.datac(!fp_functions_0_afrac_bSig_uid36_fpAddTest_b_a10_a_a13_combout),
	.datad(!fp_functions_0_areduce_nor_0_acombout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_2_a6_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_2_a6.extended_lut = "off";
defparam fp_functions_0_aMux_2_a6.lut_mask = 64'h0027002700270027;
defparam fp_functions_0_aMux_2_a6.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_afrac_bSig_uid36_fpAddTest_b_a11_a_a14(
	.dataa(!b[11]),
	.datab(!a[11]),
	.datac(!fp_functions_0_aadd_0_a1_sumout),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_afrac_bSig_uid36_fpAddTest_b_a11_a_a14_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_afrac_bSig_uid36_fpAddTest_b_a11_a_a14.extended_lut = "off";
defparam fp_functions_0_afrac_bSig_uid36_fpAddTest_b_a11_a_a14.lut_mask = 64'h5353535353535353;
defparam fp_functions_0_afrac_bSig_uid36_fpAddTest_b_a11_a_a14.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_afrac_bSig_uid36_fpAddTest_b_a12_a_a15(
	.dataa(!b[12]),
	.datab(!a[12]),
	.datac(!fp_functions_0_aadd_0_a1_sumout),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_afrac_bSig_uid36_fpAddTest_b_a12_a_a15_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_afrac_bSig_uid36_fpAddTest_b_a12_a_a15.extended_lut = "off";
defparam fp_functions_0_afrac_bSig_uid36_fpAddTest_b_a12_a_a15.lut_mask = 64'h5353535353535353;
defparam fp_functions_0_afrac_bSig_uid36_fpAddTest_b_a12_a_a15.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_2_a7(
	.dataa(!fp_functions_0_aadd_1_a11_sumout),
	.datab(!fp_functions_0_afrac_bSig_uid36_fpAddTest_b_a11_a_a14_combout),
	.datac(!fp_functions_0_afrac_bSig_uid36_fpAddTest_b_a12_a_a15_combout),
	.datad(!fp_functions_0_areduce_nor_0_acombout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_2_a7_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_2_a7.extended_lut = "off";
defparam fp_functions_0_aMux_2_a7.lut_mask = 64'h0027002700270027;
defparam fp_functions_0_aMux_2_a7.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_59_a1(
	.dataa(!fp_functions_0_aMux_2_a4_combout),
	.datab(!fp_functions_0_aMux_2_a5_combout),
	.datac(!fp_functions_0_aMux_2_a6_combout),
	.datad(!fp_functions_0_aMux_2_a7_combout),
	.datae(!fp_functions_0_aadd_1_a16_sumout),
	.dataf(!fp_functions_0_aadd_1_a21_sumout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_59_a1_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_59_a1.extended_lut = "off";
defparam fp_functions_0_aMux_59_a1.lut_mask = 64'h555533330F0F00FF;
defparam fp_functions_0_aMux_59_a1.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_2_a8(
	.dataa(!b[2]),
	.datab(!a[2]),
	.datac(!fp_functions_0_aadd_0_a1_sumout),
	.datad(!fp_functions_0_aadd_1_a11_sumout),
	.datae(!b[1]),
	.dataf(!a[1]),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_2_a8_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_2_a8.extended_lut = "off";
defparam fp_functions_0_aMux_2_a8.lut_mask = 64'h0053F0530F53FF53;
defparam fp_functions_0_aMux_2_a8.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_2_a9(
	.dataa(!fp_functions_0_aadd_1_a11_sumout),
	.datab(!b[3]),
	.datac(!a[3]),
	.datad(!fp_functions_0_aadd_0_a1_sumout),
	.datae(!b[4]),
	.dataf(!a[4]),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_2_a9_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_2_a9.extended_lut = "off";
defparam fp_functions_0_aMux_2_a9.lut_mask = 64'h220A770A225F775F;
defparam fp_functions_0_aMux_2_a9.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_afrac_bSig_uid36_fpAddTest_b_a0_a_a16(
	.dataa(!b[0]),
	.datab(!a[0]),
	.datac(!fp_functions_0_aadd_0_a1_sumout),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_afrac_bSig_uid36_fpAddTest_b_a0_a_a16_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_afrac_bSig_uid36_fpAddTest_b_a0_a_a16.extended_lut = "off";
defparam fp_functions_0_afrac_bSig_uid36_fpAddTest_b_a0_a_a16.lut_mask = 64'h5353535353535353;
defparam fp_functions_0_afrac_bSig_uid36_fpAddTest_b_a0_a_a16.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_2_a10(
	.dataa(!fp_functions_0_aadd_1_a11_sumout),
	.datab(!fp_functions_0_afrac_bSig_uid36_fpAddTest_b_a0_a_a16_combout),
	.datac(!fp_functions_0_areduce_nor_0_a0_combout),
	.datad(!fp_functions_0_areduce_nor_0_a1_combout),
	.datae(!fp_functions_0_areduce_nor_0_a2_combout),
	.dataf(!fp_functions_0_areduce_nor_0_a3_combout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_2_a10_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_2_a10.extended_lut = "off";
defparam fp_functions_0_aMux_2_a10.lut_mask = 64'h1111111111111110;
defparam fp_functions_0_aMux_2_a10.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_59_a2(
	.dataa(!fp_functions_0_aadd_1_a16_sumout),
	.datab(!fp_functions_0_aadd_1_a21_sumout),
	.datac(!fp_functions_0_aMux_2_a8_combout),
	.datad(!fp_functions_0_aMux_2_a9_combout),
	.datae(!fp_functions_0_areduce_nor_0_acombout),
	.dataf(!fp_functions_0_aMux_2_a10_combout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_59_a2_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_59_a2.extended_lut = "off";
defparam fp_functions_0_aMux_59_a2.lut_mask = 64'h0000021344444657;
defparam fp_functions_0_aMux_59_a2.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_afrac_bSig_uid36_fpAddTest_b_a21_a_a17(
	.dataa(!b[21]),
	.datab(!a[21]),
	.datac(!fp_functions_0_aadd_0_a1_sumout),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_afrac_bSig_uid36_fpAddTest_b_a21_a_a17_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_afrac_bSig_uid36_fpAddTest_b_a21_a_a17.extended_lut = "off";
defparam fp_functions_0_afrac_bSig_uid36_fpAddTest_b_a21_a_a17.lut_mask = 64'h5353535353535353;
defparam fp_functions_0_afrac_bSig_uid36_fpAddTest_b_a21_a_a17.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_2_a11(
	.dataa(!fp_functions_0_aadd_1_a11_sumout),
	.datab(!fp_functions_0_areduce_nor_0_a0_combout),
	.datac(!fp_functions_0_areduce_nor_0_a1_combout),
	.datad(!fp_functions_0_areduce_nor_0_a2_combout),
	.datae(!fp_functions_0_areduce_nor_0_a3_combout),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_2_a11_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_2_a11.extended_lut = "off";
defparam fp_functions_0_aMux_2_a11.lut_mask = 64'hAAAAAAA8AAAAAAA8;
defparam fp_functions_0_aMux_2_a11.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_afrac_bSig_uid36_fpAddTest_b_a22_a_a18(
	.dataa(!b[22]),
	.datab(!a[22]),
	.datac(!fp_functions_0_aadd_0_a1_sumout),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_afrac_bSig_uid36_fpAddTest_b_a22_a_a18_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_afrac_bSig_uid36_fpAddTest_b_a22_a_a18.extended_lut = "off";
defparam fp_functions_0_afrac_bSig_uid36_fpAddTest_b_a22_a_a18.lut_mask = 64'h5353535353535353;
defparam fp_functions_0_afrac_bSig_uid36_fpAddTest_b_a22_a_a18.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_2_a12(
	.dataa(!fp_functions_0_aadd_1_a11_sumout),
	.datab(!fp_functions_0_afrac_bSig_uid36_fpAddTest_b_a22_a_a18_combout),
	.datac(!fp_functions_0_areduce_nor_0_a0_combout),
	.datad(!fp_functions_0_areduce_nor_0_a1_combout),
	.datae(!fp_functions_0_areduce_nor_0_a2_combout),
	.dataf(!fp_functions_0_areduce_nor_0_a3_combout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_2_a12_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_2_a12.extended_lut = "off";
defparam fp_functions_0_aMux_2_a12.lut_mask = 64'h1111111111111110;
defparam fp_functions_0_aMux_2_a12.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_59_a3(
	.dataa(!fp_functions_0_afrac_bSig_uid36_fpAddTest_b_a21_a_a17_combout),
	.datab(!fp_functions_0_aadd_1_a16_sumout),
	.datac(!fp_functions_0_aadd_1_a21_sumout),
	.datad(!fp_functions_0_aadd_1_a1_sumout),
	.datae(!fp_functions_0_aMux_2_a11_combout),
	.dataf(!fp_functions_0_aMux_2_a12_combout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_59_a3_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_59_a3.extended_lut = "off";
defparam fp_functions_0_aMux_59_a3.lut_mask = 64'h0000007000C000F0;
defparam fp_functions_0_aMux_59_a3.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai1783_a0(
	.dataa(!fp_functions_0_aadd_1_a1_sumout),
	.datab(!fp_functions_0_aadd_1_a6_sumout),
	.datac(!fp_functions_0_aMux_59_a0_combout),
	.datad(!fp_functions_0_aMux_59_a1_combout),
	.datae(!fp_functions_0_aMux_59_a2_combout),
	.dataf(!fp_functions_0_aMux_59_a3_combout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai1783_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai1783_a0.extended_lut = "off";
defparam fp_functions_0_ai1783_a0.lut_mask = 64'h02468ACE3377BBFF;
defparam fp_functions_0_ai1783_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a28_a_a0(
	.dataa(!areset),
	.datab(!fp_functions_0_aadd_1_a26_sumout),
	.datac(!fp_functions_0_aadd_3_a1_sumout),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a28_a_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a28_a_a0.extended_lut = "off";
defparam fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a28_a_a0.lut_mask = 64'hF7F7F7F7F7F7F7F7;
defparam fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a28_a_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_2_a13(
	.dataa(!fp_functions_0_aadd_1_a11_sumout),
	.datab(!fp_functions_0_afrac_bSig_uid36_fpAddTest_b_a21_a_a17_combout),
	.datac(!fp_functions_0_afrac_bSig_uid36_fpAddTest_b_a22_a_a18_combout),
	.datad(!fp_functions_0_areduce_nor_0_acombout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_2_a13_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_2_a13.extended_lut = "off";
defparam fp_functions_0_aMux_2_a13.lut_mask = 64'h0027002700270027;
defparam fp_functions_0_aMux_2_a13.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_57_a0(
	.dataa(!fp_functions_0_aMux_2_a1_combout),
	.datab(!fp_functions_0_aMux_2_a2_combout),
	.datac(!fp_functions_0_aMux_2_a3_combout),
	.datad(!fp_functions_0_aMux_2_a13_combout),
	.datae(!fp_functions_0_aadd_1_a16_sumout),
	.dataf(!fp_functions_0_aadd_1_a21_sumout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_57_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_57_a0.extended_lut = "off";
defparam fp_functions_0_aMux_57_a0.lut_mask = 64'h555533330F0F00FF;
defparam fp_functions_0_aMux_57_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_57_a1(
	.dataa(!fp_functions_0_aMux_2_a5_combout),
	.datab(!fp_functions_0_aMux_2_a6_combout),
	.datac(!fp_functions_0_aMux_2_a7_combout),
	.datad(!fp_functions_0_aMux_2_a0_combout),
	.datae(!fp_functions_0_aadd_1_a16_sumout),
	.dataf(!fp_functions_0_aadd_1_a21_sumout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_57_a1_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_57_a1.extended_lut = "off";
defparam fp_functions_0_aMux_57_a1.lut_mask = 64'h555533330F0F00FF;
defparam fp_functions_0_aMux_57_a1.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_65_a0(
	.dataa(!fp_functions_0_aadd_1_a1_sumout),
	.datab(!fp_functions_0_aMux_57_a0_combout),
	.datac(!fp_functions_0_aMux_57_a1_combout),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_65_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_65_a0.extended_lut = "off";
defparam fp_functions_0_aMux_65_a0.lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam fp_functions_0_aMux_65_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_2_a14(
	.dataa(!fp_functions_0_aMux_2_a8_combout),
	.datab(!fp_functions_0_areduce_nor_0_acombout),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_2_a14_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_2_a14.extended_lut = "off";
defparam fp_functions_0_aMux_2_a14.lut_mask = 64'h1111111111111111;
defparam fp_functions_0_aMux_2_a14.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_2_a15(
	.dataa(!fp_functions_0_aMux_2_a9_combout),
	.datab(!fp_functions_0_areduce_nor_0_acombout),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_2_a15_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_2_a15.extended_lut = "off";
defparam fp_functions_0_aMux_2_a15.lut_mask = 64'h1111111111111111;
defparam fp_functions_0_aMux_2_a15.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_57_a2(
	.dataa(!fp_functions_0_aMux_2_a10_combout),
	.datab(!fp_functions_0_aadd_1_a16_sumout),
	.datac(!fp_functions_0_aadd_1_a21_sumout),
	.datad(!fp_functions_0_aMux_2_a4_combout),
	.datae(!fp_functions_0_aMux_2_a14_combout),
	.dataf(!fp_functions_0_aMux_2_a15_combout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_57_a2_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_57_a2.extended_lut = "off";
defparam fp_functions_0_aMux_57_a2.lut_mask = 64'h404370734C4F7C7F;
defparam fp_functions_0_aMux_57_a2.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_49_a0(
	.dataa(!fp_functions_0_aadd_1_a16_sumout),
	.datab(!fp_functions_0_aadd_1_a21_sumout),
	.datac(!fp_functions_0_aadd_1_a1_sumout),
	.datad(!fp_functions_0_aMux_2_a11_combout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_49_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_49_a0.extended_lut = "off";
defparam fp_functions_0_aMux_49_a0.lut_mask = 64'h0080008000800080;
defparam fp_functions_0_aMux_49_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai1734_a0(
	.dataa(!fp_functions_0_aadd_1_a1_sumout),
	.datab(!fp_functions_0_aadd_1_a26_sumout),
	.datac(!fp_functions_0_aMux_57_a2_combout),
	.datad(!fp_functions_0_aMux_49_a0_combout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai1734_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai1734_a0.extended_lut = "off";
defparam fp_functions_0_ai1734_a0.lut_mask = 64'h0437043704370437;
defparam fp_functions_0_ai1734_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai1734_a1(
	.dataa(!fp_functions_0_aadd_1_a6_sumout),
	.datab(!fp_functions_0_aadd_1_a26_sumout),
	.datac(!fp_functions_0_aMux_65_a0_combout),
	.datad(!fp_functions_0_ai1734_a0_combout),
	.datae(!fp_functions_0_aadd_3_a1_sumout),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai1734_a1_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai1734_a1.extended_lut = "off";
defparam fp_functions_0_ai1734_a1.lut_mask = 64'h000004AE000004AE;
defparam fp_functions_0_ai1734_a1.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai1734_a2(
	.dataa(!fp_functions_0_aadd_1_a6_sumout),
	.datab(!fp_functions_0_aadd_1_a26_sumout),
	.datac(!fp_functions_0_aMux_65_a0_combout),
	.datad(!fp_functions_0_ai1734_a0_combout),
	.datae(!fp_functions_0_aadd_3_a1_sumout),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai1734_a2_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai1734_a2.extended_lut = "off";
defparam fp_functions_0_ai1734_a2.lut_mask = 64'h0000025700000257;
defparam fp_functions_0_ai1734_a2.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_2_a16(
	.dataa(!fp_functions_0_aadd_1_a11_sumout),
	.datab(!fp_functions_0_afrac_bSig_uid36_fpAddTest_b_a16_a_a3_combout),
	.datac(!fp_functions_0_afrac_bSig_uid36_fpAddTest_b_a17_a_a4_combout),
	.datad(!fp_functions_0_areduce_nor_0_acombout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_2_a16_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_2_a16.extended_lut = "off";
defparam fp_functions_0_aMux_2_a16.lut_mask = 64'h0027002700270027;
defparam fp_functions_0_aMux_2_a16.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_2_a17(
	.dataa(!fp_functions_0_aadd_1_a11_sumout),
	.datab(!b[20]),
	.datac(!a[20]),
	.datad(!fp_functions_0_aadd_0_a1_sumout),
	.datae(!b[21]),
	.dataf(!a[21]),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_2_a17_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_2_a17.extended_lut = "off";
defparam fp_functions_0_aMux_2_a17.lut_mask = 64'h220A770A225F775F;
defparam fp_functions_0_aMux_2_a17.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_2_a18(
	.dataa(!fp_functions_0_aMux_2_a17_combout),
	.datab(!fp_functions_0_areduce_nor_0_acombout),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_2_a18_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_2_a18.extended_lut = "off";
defparam fp_functions_0_aMux_2_a18.lut_mask = 64'h1111111111111111;
defparam fp_functions_0_aMux_2_a18.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_2_a19(
	.dataa(!fp_functions_0_aadd_1_a11_sumout),
	.datab(!fp_functions_0_afrac_bSig_uid36_fpAddTest_b_a18_a_a5_combout),
	.datac(!fp_functions_0_afrac_bSig_uid36_fpAddTest_b_a19_a_a6_combout),
	.datad(!fp_functions_0_areduce_nor_0_acombout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_2_a19_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_2_a19.extended_lut = "off";
defparam fp_functions_0_aMux_2_a19.lut_mask = 64'h0027002700270027;
defparam fp_functions_0_aMux_2_a19.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_2_a20(
	.dataa(!fp_functions_0_aadd_1_a11_sumout),
	.datab(!fp_functions_0_afrac_bSig_uid36_fpAddTest_b_a22_a_a18_combout),
	.datac(!fp_functions_0_areduce_nor_0_a0_combout),
	.datad(!fp_functions_0_areduce_nor_0_a1_combout),
	.datae(!fp_functions_0_areduce_nor_0_a2_combout),
	.dataf(!fp_functions_0_areduce_nor_0_a3_combout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_2_a20_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_2_a20.extended_lut = "off";
defparam fp_functions_0_aMux_2_a20.lut_mask = 64'h888888888888888F;
defparam fp_functions_0_aMux_2_a20.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_60_a0(
	.dataa(!fp_functions_0_aMux_2_a16_combout),
	.datab(!fp_functions_0_aMux_2_a18_combout),
	.datac(!fp_functions_0_aMux_2_a19_combout),
	.datad(!fp_functions_0_aMux_2_a20_combout),
	.datae(!fp_functions_0_aadd_1_a21_sumout),
	.dataf(!fp_functions_0_aadd_1_a16_sumout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_60_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_60_a0.extended_lut = "off";
defparam fp_functions_0_aMux_60_a0.lut_mask = 64'h555533330F0FFF00;
defparam fp_functions_0_aMux_60_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_2_a21(
	.dataa(!fp_functions_0_aadd_1_a11_sumout),
	.datab(!fp_functions_0_afrac_bSig_uid36_fpAddTest_b_a8_a_a11_combout),
	.datac(!fp_functions_0_afrac_bSig_uid36_fpAddTest_b_a9_a_a12_combout),
	.datad(!fp_functions_0_areduce_nor_0_acombout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_2_a21_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_2_a21.extended_lut = "off";
defparam fp_functions_0_aMux_2_a21.lut_mask = 64'h0027002700270027;
defparam fp_functions_0_aMux_2_a21.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_2_a22(
	.dataa(!fp_functions_0_aadd_1_a11_sumout),
	.datab(!fp_functions_0_afrac_bSig_uid36_fpAddTest_b_a10_a_a13_combout),
	.datac(!fp_functions_0_afrac_bSig_uid36_fpAddTest_b_a11_a_a14_combout),
	.datad(!fp_functions_0_areduce_nor_0_acombout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_2_a22_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_2_a22.extended_lut = "off";
defparam fp_functions_0_aMux_2_a22.lut_mask = 64'h0027002700270027;
defparam fp_functions_0_aMux_2_a22.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_2_a23(
	.dataa(!fp_functions_0_aadd_1_a11_sumout),
	.datab(!fp_functions_0_afrac_bSig_uid36_fpAddTest_b_a12_a_a15_combout),
	.datac(!fp_functions_0_afrac_bSig_uid36_fpAddTest_b_a13_a_a0_combout),
	.datad(!fp_functions_0_areduce_nor_0_acombout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_2_a23_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_2_a23.extended_lut = "off";
defparam fp_functions_0_aMux_2_a23.lut_mask = 64'h0027002700270027;
defparam fp_functions_0_aMux_2_a23.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_2_a24(
	.dataa(!fp_functions_0_aadd_1_a11_sumout),
	.datab(!fp_functions_0_afrac_bSig_uid36_fpAddTest_b_a14_a_a1_combout),
	.datac(!fp_functions_0_afrac_bSig_uid36_fpAddTest_b_a15_a_a2_combout),
	.datad(!fp_functions_0_areduce_nor_0_acombout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_2_a24_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_2_a24.extended_lut = "off";
defparam fp_functions_0_aMux_2_a24.lut_mask = 64'h0027002700270027;
defparam fp_functions_0_aMux_2_a24.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_60_a1(
	.dataa(!fp_functions_0_aMux_2_a21_combout),
	.datab(!fp_functions_0_aMux_2_a22_combout),
	.datac(!fp_functions_0_aMux_2_a23_combout),
	.datad(!fp_functions_0_aMux_2_a24_combout),
	.datae(!fp_functions_0_aadd_1_a16_sumout),
	.dataf(!fp_functions_0_aadd_1_a21_sumout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_60_a1_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_60_a1.extended_lut = "off";
defparam fp_functions_0_aMux_60_a1.lut_mask = 64'h555533330F0F00FF;
defparam fp_functions_0_aMux_60_a1.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_23_a0(
	.dataa(!b[1]),
	.datab(!a[1]),
	.datac(!fp_functions_0_aadd_0_a1_sumout),
	.datad(!fp_functions_0_aadd_1_a11_sumout),
	.datae(!fp_functions_0_afrac_bSig_uid36_fpAddTest_b_a0_a_a16_combout),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_23_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_23_a0.extended_lut = "off";
defparam fp_functions_0_aMux_23_a0.lut_mask = 64'h0053FF530053FF53;
defparam fp_functions_0_aMux_23_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_2_a25(
	.dataa(!fp_functions_0_aMux_23_a0_combout),
	.datab(!fp_functions_0_areduce_nor_0_acombout),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_2_a25_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_2_a25.extended_lut = "off";
defparam fp_functions_0_aMux_2_a25.lut_mask = 64'h1111111111111111;
defparam fp_functions_0_aMux_2_a25.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_2_a26(
	.dataa(!fp_functions_0_aadd_1_a11_sumout),
	.datab(!b[4]),
	.datac(!a[4]),
	.datad(!fp_functions_0_aadd_0_a1_sumout),
	.datae(!b[5]),
	.dataf(!a[5]),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_2_a26_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_2_a26.extended_lut = "off";
defparam fp_functions_0_aMux_2_a26.lut_mask = 64'h220A770A225F775F;
defparam fp_functions_0_aMux_2_a26.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_2_a27(
	.dataa(!fp_functions_0_aMux_2_a26_combout),
	.datab(!fp_functions_0_areduce_nor_0_acombout),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_2_a27_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_2_a27.extended_lut = "off";
defparam fp_functions_0_aMux_2_a27.lut_mask = 64'h1111111111111111;
defparam fp_functions_0_aMux_2_a27.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_23_a1(
	.dataa(!b[2]),
	.datab(!a[2]),
	.datac(!fp_functions_0_aadd_0_a1_sumout),
	.datad(!fp_functions_0_aadd_1_a11_sumout),
	.datae(!b[3]),
	.dataf(!a[3]),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_23_a1_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_23_a1.extended_lut = "off";
defparam fp_functions_0_aMux_23_a1.lut_mask = 64'h530053F0530F53FF;
defparam fp_functions_0_aMux_23_a1.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_2_a28(
	.dataa(!fp_functions_0_aMux_23_a1_combout),
	.datab(!fp_functions_0_areduce_nor_0_acombout),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_2_a28_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_2_a28.extended_lut = "off";
defparam fp_functions_0_aMux_2_a28.lut_mask = 64'h1111111111111111;
defparam fp_functions_0_aMux_2_a28.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_2_a29(
	.dataa(!fp_functions_0_aadd_1_a11_sumout),
	.datab(!fp_functions_0_afrac_bSig_uid36_fpAddTest_b_a7_a_a10_combout),
	.datac(!fp_functions_0_afrac_bSig_uid36_fpAddTest_b_a6_a_a9_combout),
	.datad(!fp_functions_0_areduce_nor_0_acombout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_2_a29_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_2_a29.extended_lut = "off";
defparam fp_functions_0_aMux_2_a29.lut_mask = 64'h001B001B001B001B;
defparam fp_functions_0_aMux_2_a29.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_60_a2(
	.dataa(!fp_functions_0_aMux_2_a25_combout),
	.datab(!fp_functions_0_aMux_2_a27_combout),
	.datac(!fp_functions_0_aMux_2_a28_combout),
	.datad(!fp_functions_0_aMux_2_a29_combout),
	.datae(!fp_functions_0_aadd_1_a21_sumout),
	.dataf(!fp_functions_0_aadd_1_a16_sumout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_60_a2_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_60_a2.extended_lut = "off";
defparam fp_functions_0_aMux_60_a2.lut_mask = 64'h555533330F0F00FF;
defparam fp_functions_0_aMux_60_a2.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai1783_a1(
	.dataa(!fp_functions_0_aadd_1_a1_sumout),
	.datab(!fp_functions_0_aadd_1_a26_sumout),
	.datac(!fp_functions_0_aMux_60_a0_combout),
	.datad(!fp_functions_0_aMux_60_a1_combout),
	.datae(!fp_functions_0_aMux_60_a2_combout),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai1783_a1_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai1783_a1.extended_lut = "off";
defparam fp_functions_0_ai1783_a1.lut_mask = 64'h0123456701234567;
defparam fp_functions_0_ai1783_a1.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a2_a_a1(
	.dataa(!areset),
	.datab(!fp_functions_0_aadd_1_a6_sumout),
	.datac(!fp_functions_0_aadd_1_a26_sumout),
	.datad(!fp_functions_0_aadd_3_a1_sumout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a2_a_a1_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a2_a_a1.extended_lut = "off";
defparam fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a2_a_a1.lut_mask = 64'hFFD7FFD7FFD7FFD7;
defparam fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a2_a_a1.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai1783_a2(
	.dataa(!fp_functions_0_aadd_1_a1_sumout),
	.datab(!fp_functions_0_aadd_1_a26_sumout),
	.datac(!fp_functions_0_aMux_60_a0_combout),
	.datad(!fp_functions_0_aMux_60_a1_combout),
	.datae(!fp_functions_0_aMux_60_a2_combout),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai1783_a2_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai1783_a2.extended_lut = "off";
defparam fp_functions_0_ai1783_a2.lut_mask = 64'h02468ACE02468ACE;
defparam fp_functions_0_ai1783_a2.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_57_a3(
	.dataa(!fp_functions_0_aMux_2_a7_combout),
	.datab(!fp_functions_0_aMux_2_a0_combout),
	.datac(!fp_functions_0_aMux_2_a1_combout),
	.datad(!fp_functions_0_aMux_2_a2_combout),
	.datae(!fp_functions_0_aadd_1_a16_sumout),
	.dataf(!fp_functions_0_aadd_1_a21_sumout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_57_a3_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_57_a3.extended_lut = "off";
defparam fp_functions_0_aMux_57_a3.lut_mask = 64'h555533330F0F00FF;
defparam fp_functions_0_aMux_57_a3.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_57_a4(
	.dataa(!fp_functions_0_aMux_2_a15_combout),
	.datab(!fp_functions_0_aMux_2_a4_combout),
	.datac(!fp_functions_0_aMux_2_a5_combout),
	.datad(!fp_functions_0_aMux_2_a6_combout),
	.datae(!fp_functions_0_aadd_1_a16_sumout),
	.dataf(!fp_functions_0_aadd_1_a21_sumout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_57_a4_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_57_a4.extended_lut = "off";
defparam fp_functions_0_aMux_57_a4.lut_mask = 64'h555533330F0F00FF;
defparam fp_functions_0_aMux_57_a4.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_61_a0(
	.dataa(!fp_functions_0_aadd_1_a16_sumout),
	.datab(!fp_functions_0_aadd_1_a21_sumout),
	.datac(!fp_functions_0_aadd_1_a1_sumout),
	.datad(!fp_functions_0_aMux_2_a11_combout),
	.datae(!fp_functions_0_aMux_2_a3_combout),
	.dataf(!fp_functions_0_aMux_2_a13_combout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_61_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_61_a0.extended_lut = "off";
defparam fp_functions_0_aMux_61_a0.lut_mask = 64'h0002080A04060C0E;
defparam fp_functions_0_aMux_61_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_77_a0(
	.dataa(!fp_functions_0_aadd_1_a16_sumout),
	.datab(!fp_functions_0_aadd_1_a21_sumout),
	.datac(!fp_functions_0_aMux_2_a8_combout),
	.datad(!fp_functions_0_aadd_1_a1_sumout),
	.datae(!fp_functions_0_areduce_nor_0_acombout),
	.dataf(!fp_functions_0_aMux_2_a10_combout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_77_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_77_a0.extended_lut = "off";
defparam fp_functions_0_aMux_77_a0.lut_mask = 64'h0000010022002300;
defparam fp_functions_0_aMux_77_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai1783_a3(
	.dataa(!fp_functions_0_aadd_1_a1_sumout),
	.datab(!fp_functions_0_aadd_1_a26_sumout),
	.datac(!fp_functions_0_aMux_57_a3_combout),
	.datad(!fp_functions_0_aMux_57_a4_combout),
	.datae(!fp_functions_0_aMux_61_a0_combout),
	.dataf(!fp_functions_0_aMux_77_a0_combout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai1783_a3_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai1783_a3.extended_lut = "off";
defparam fp_functions_0_ai1783_a3.lut_mask = 64'h02463377CECEFFFF;
defparam fp_functions_0_ai1783_a3.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_60_a3(
	.dataa(!fp_functions_0_aMux_2_a23_combout),
	.datab(!fp_functions_0_aMux_2_a24_combout),
	.datac(!fp_functions_0_aMux_2_a16_combout),
	.datad(!fp_functions_0_aMux_2_a19_combout),
	.datae(!fp_functions_0_aadd_1_a16_sumout),
	.dataf(!fp_functions_0_aadd_1_a21_sumout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_60_a3_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_60_a3.extended_lut = "off";
defparam fp_functions_0_aMux_60_a3.lut_mask = 64'h555533330F0F00FF;
defparam fp_functions_0_aMux_60_a3.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_60_a4(
	.dataa(!fp_functions_0_aMux_2_a27_combout),
	.datab(!fp_functions_0_aMux_2_a29_combout),
	.datac(!fp_functions_0_aMux_2_a21_combout),
	.datad(!fp_functions_0_aMux_2_a22_combout),
	.datae(!fp_functions_0_aadd_1_a16_sumout),
	.dataf(!fp_functions_0_aadd_1_a21_sumout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_60_a4_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_60_a4.extended_lut = "off";
defparam fp_functions_0_aMux_60_a4.lut_mask = 64'h555533330F0F00FF;
defparam fp_functions_0_aMux_60_a4.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_76_a0(
	.dataa(!fp_functions_0_aadd_1_a16_sumout),
	.datab(!fp_functions_0_aadd_1_a21_sumout),
	.datac(!fp_functions_0_aMux_23_a0_combout),
	.datad(!fp_functions_0_aMux_23_a1_combout),
	.datae(!fp_functions_0_aadd_1_a1_sumout),
	.dataf(!fp_functions_0_areduce_nor_0_acombout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_76_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_76_a0.extended_lut = "off";
defparam fp_functions_0_aMux_76_a0.lut_mask = 64'h0000000002130000;
defparam fp_functions_0_aMux_76_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_60_a5(
	.dataa(!fp_functions_0_aadd_1_a16_sumout),
	.datab(!fp_functions_0_aadd_1_a21_sumout),
	.datac(!fp_functions_0_aMux_2_a17_combout),
	.datad(!fp_functions_0_aadd_1_a1_sumout),
	.datae(!fp_functions_0_areduce_nor_0_acombout),
	.dataf(!fp_functions_0_aMux_2_a20_combout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_60_a5_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_60_a5.extended_lut = "off";
defparam fp_functions_0_aMux_60_a5.lut_mask = 64'h0044004C00000008;
defparam fp_functions_0_aMux_60_a5.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai1783_a4(
	.dataa(!fp_functions_0_aadd_1_a1_sumout),
	.datab(!fp_functions_0_aadd_1_a6_sumout),
	.datac(!fp_functions_0_aMux_60_a3_combout),
	.datad(!fp_functions_0_aMux_60_a4_combout),
	.datae(!fp_functions_0_aMux_76_a0_combout),
	.dataf(!fp_functions_0_aMux_60_a5_combout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai1783_a4_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai1783_a4.extended_lut = "off";
defparam fp_functions_0_ai1783_a4.lut_mask = 64'h0246CECE3377FFFF;
defparam fp_functions_0_ai1783_a4.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai1783_a5(
	.dataa(!fp_functions_0_aadd_1_a1_sumout),
	.datab(!fp_functions_0_aadd_1_a6_sumout),
	.datac(!fp_functions_0_aMux_57_a3_combout),
	.datad(!fp_functions_0_aMux_57_a4_combout),
	.datae(!fp_functions_0_aMux_61_a0_combout),
	.dataf(!fp_functions_0_aMux_77_a0_combout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai1783_a5_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai1783_a5.extended_lut = "off";
defparam fp_functions_0_ai1783_a5.lut_mask = 64'h02463377CECEFFFF;
defparam fp_functions_0_ai1783_a5.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_58_a0(
	.dataa(!fp_functions_0_aMux_2_a22_combout),
	.datab(!fp_functions_0_aMux_2_a23_combout),
	.datac(!fp_functions_0_aMux_2_a24_combout),
	.datad(!fp_functions_0_aMux_2_a16_combout),
	.datae(!fp_functions_0_aadd_1_a16_sumout),
	.dataf(!fp_functions_0_aadd_1_a21_sumout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_58_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_58_a0.extended_lut = "off";
defparam fp_functions_0_aMux_58_a0.lut_mask = 64'h555533330F0F00FF;
defparam fp_functions_0_aMux_58_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_58_a1(
	.dataa(!fp_functions_0_aMux_2_a28_combout),
	.datab(!fp_functions_0_aMux_2_a27_combout),
	.datac(!fp_functions_0_aMux_2_a29_combout),
	.datad(!fp_functions_0_aMux_2_a21_combout),
	.datae(!fp_functions_0_aadd_1_a16_sumout),
	.dataf(!fp_functions_0_aadd_1_a21_sumout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_58_a1_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_58_a1.extended_lut = "off";
defparam fp_functions_0_aMux_58_a1.lut_mask = 64'h555533330F0F00FF;
defparam fp_functions_0_aMux_58_a1.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_78_a0(
	.dataa(!fp_functions_0_aadd_1_a16_sumout),
	.datab(!fp_functions_0_aadd_1_a21_sumout),
	.datac(!fp_functions_0_aMux_23_a0_combout),
	.datad(!fp_functions_0_aadd_1_a1_sumout),
	.datae(!fp_functions_0_areduce_nor_0_acombout),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_78_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_78_a0.extended_lut = "off";
defparam fp_functions_0_aMux_78_a0.lut_mask = 64'h0000010000000100;
defparam fp_functions_0_aMux_78_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_62_a0(
	.dataa(!fp_functions_0_aadd_1_a16_sumout),
	.datab(!fp_functions_0_aadd_1_a21_sumout),
	.datac(!fp_functions_0_aadd_1_a1_sumout),
	.datad(!fp_functions_0_aMux_2_a19_combout),
	.datae(!fp_functions_0_aMux_2_a20_combout),
	.dataf(!fp_functions_0_aMux_2_a18_combout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_62_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_62_a0.extended_lut = "off";
defparam fp_functions_0_aMux_62_a0.lut_mask = 64'h020A0008060E040C;
defparam fp_functions_0_aMux_62_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai1783_a6(
	.dataa(!fp_functions_0_aadd_1_a1_sumout),
	.datab(!fp_functions_0_aadd_1_a6_sumout),
	.datac(!fp_functions_0_aMux_58_a0_combout),
	.datad(!fp_functions_0_aMux_58_a1_combout),
	.datae(!fp_functions_0_aMux_78_a0_combout),
	.dataf(!fp_functions_0_aMux_62_a0_combout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai1783_a6_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai1783_a6.extended_lut = "off";
defparam fp_functions_0_ai1783_a6.lut_mask = 64'h0246CECE3377FFFF;
defparam fp_functions_0_ai1783_a6.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai1783_a7(
	.dataa(!fp_functions_0_aadd_1_a1_sumout),
	.datab(!fp_functions_0_aadd_1_a6_sumout),
	.datac(!fp_functions_0_aMux_60_a0_combout),
	.datad(!fp_functions_0_aMux_60_a1_combout),
	.datae(!fp_functions_0_aMux_60_a2_combout),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai1783_a7_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai1783_a7.extended_lut = "off";
defparam fp_functions_0_ai1783_a7.lut_mask = 64'h0123456701234567;
defparam fp_functions_0_ai1783_a7.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_59_a4(
	.dataa(!fp_functions_0_aMux_2_a11_combout),
	.datab(!fp_functions_0_aadd_1_a16_sumout),
	.datac(!fp_functions_0_aadd_1_a21_sumout),
	.datad(!fp_functions_0_aMux_2_a3_combout),
	.datae(!fp_functions_0_aMux_2_a13_combout),
	.dataf(!fp_functions_0_aMux_2_a2_combout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_59_a4_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_59_a4.extended_lut = "off";
defparam fp_functions_0_aMux_59_a4.lut_mask = 64'h01310D3DC1F1CDFD;
defparam fp_functions_0_aMux_59_a4.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_59_a5(
	.dataa(!fp_functions_0_aMux_2_a6_combout),
	.datab(!fp_functions_0_aMux_2_a7_combout),
	.datac(!fp_functions_0_aMux_2_a0_combout),
	.datad(!fp_functions_0_aMux_2_a1_combout),
	.datae(!fp_functions_0_aadd_1_a16_sumout),
	.dataf(!fp_functions_0_aadd_1_a21_sumout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_59_a5_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_59_a5.extended_lut = "off";
defparam fp_functions_0_aMux_59_a5.lut_mask = 64'h555533330F0F00FF;
defparam fp_functions_0_aMux_59_a5.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_59_a6(
	.dataa(!fp_functions_0_aMux_2_a14_combout),
	.datab(!fp_functions_0_aMux_2_a15_combout),
	.datac(!fp_functions_0_aMux_2_a4_combout),
	.datad(!fp_functions_0_aMux_2_a5_combout),
	.datae(!fp_functions_0_aadd_1_a16_sumout),
	.dataf(!fp_functions_0_aadd_1_a21_sumout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_59_a6_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_59_a6.extended_lut = "off";
defparam fp_functions_0_aMux_59_a6.lut_mask = 64'h555533330F0F00FF;
defparam fp_functions_0_aMux_59_a6.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_79_a0(
	.dataa(!fp_functions_0_aadd_1_a16_sumout),
	.datab(!fp_functions_0_aadd_1_a21_sumout),
	.datac(!fp_functions_0_aadd_1_a1_sumout),
	.datad(!fp_functions_0_aMux_2_a10_combout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_79_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_79_a0.extended_lut = "off";
defparam fp_functions_0_aMux_79_a0.lut_mask = 64'h0010001000100010;
defparam fp_functions_0_aMux_79_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai1783_a8(
	.dataa(!fp_functions_0_aadd_1_a1_sumout),
	.datab(!fp_functions_0_aadd_1_a6_sumout),
	.datac(!fp_functions_0_aMux_59_a4_combout),
	.datad(!fp_functions_0_aMux_59_a5_combout),
	.datae(!fp_functions_0_aMux_59_a6_combout),
	.dataf(!fp_functions_0_aMux_79_a0_combout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai1783_a8_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai1783_a8.extended_lut = "off";
defparam fp_functions_0_ai1783_a8.lut_mask = 64'h01234567CDEFCDEF;
defparam fp_functions_0_ai1783_a8.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_57_a5(
	.dataa(!fp_functions_0_aadd_1_a16_sumout),
	.datab(!fp_functions_0_aadd_1_a21_sumout),
	.datac(!fp_functions_0_aadd_1_a1_sumout),
	.datad(!fp_functions_0_aMux_2_a11_combout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_57_a5_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_57_a5.extended_lut = "off";
defparam fp_functions_0_aMux_57_a5.lut_mask = 64'h0008000800080008;
defparam fp_functions_0_aMux_57_a5.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai1783_a9(
	.dataa(!fp_functions_0_aadd_1_a1_sumout),
	.datab(!fp_functions_0_aadd_1_a26_sumout),
	.datac(!fp_functions_0_aMux_57_a0_combout),
	.datad(!fp_functions_0_aMux_57_a1_combout),
	.datae(!fp_functions_0_aMux_57_a5_combout),
	.dataf(!fp_functions_0_aMux_57_a2_combout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai1783_a9_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai1783_a9.extended_lut = "off";
defparam fp_functions_0_ai1783_a9.lut_mask = 64'h024633778ACEBBFF;
defparam fp_functions_0_ai1783_a9.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_58_a2(
	.dataa(!fp_functions_0_aMux_2_a24_combout),
	.datab(!fp_functions_0_aMux_2_a16_combout),
	.datac(!fp_functions_0_aMux_2_a19_combout),
	.datad(!fp_functions_0_aMux_2_a18_combout),
	.datae(!fp_functions_0_aadd_1_a16_sumout),
	.dataf(!fp_functions_0_aadd_1_a21_sumout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_58_a2_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_58_a2.extended_lut = "off";
defparam fp_functions_0_aMux_58_a2.lut_mask = 64'h555533330F0F00FF;
defparam fp_functions_0_aMux_58_a2.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_58_a3(
	.dataa(!fp_functions_0_aMux_2_a29_combout),
	.datab(!fp_functions_0_aMux_2_a21_combout),
	.datac(!fp_functions_0_aMux_2_a22_combout),
	.datad(!fp_functions_0_aMux_2_a23_combout),
	.datae(!fp_functions_0_aadd_1_a16_sumout),
	.dataf(!fp_functions_0_aadd_1_a21_sumout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_58_a3_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_58_a3.extended_lut = "off";
defparam fp_functions_0_aMux_58_a3.lut_mask = 64'h555533330F0F00FF;
defparam fp_functions_0_aMux_58_a3.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_58_a4(
	.dataa(!fp_functions_0_aadd_1_a16_sumout),
	.datab(!fp_functions_0_aadd_1_a21_sumout),
	.datac(!fp_functions_0_aadd_1_a1_sumout),
	.datad(!fp_functions_0_aMux_2_a20_combout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_58_a4_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_58_a4.extended_lut = "off";
defparam fp_functions_0_aMux_58_a4.lut_mask = 64'h0800080008000800;
defparam fp_functions_0_aMux_58_a4.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai1783_a10(
	.dataa(!fp_functions_0_aadd_1_a16_sumout),
	.datab(!fp_functions_0_aadd_1_a21_sumout),
	.datac(!fp_functions_0_aadd_1_a1_sumout),
	.datad(!fp_functions_0_aMux_2_a25_combout),
	.datae(!fp_functions_0_aMux_2_a28_combout),
	.dataf(!fp_functions_0_aMux_2_a27_combout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai1783_a10_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai1783_a10.extended_lut = "off";
defparam fp_functions_0_ai1783_a10.lut_mask = 64'h0040206010503070;
defparam fp_functions_0_ai1783_a10.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai1783_a11(
	.dataa(!fp_functions_0_aadd_1_a1_sumout),
	.datab(!fp_functions_0_aadd_1_a26_sumout),
	.datac(!fp_functions_0_aMux_58_a2_combout),
	.datad(!fp_functions_0_aMux_58_a3_combout),
	.datae(!fp_functions_0_aMux_58_a4_combout),
	.dataf(!fp_functions_0_ai1783_a10_combout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai1783_a11_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai1783_a11.extended_lut = "off";
defparam fp_functions_0_ai1783_a11.lut_mask = 64'h02463377CECEFFFF;
defparam fp_functions_0_ai1783_a11.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai1783_a12(
	.dataa(!fp_functions_0_aadd_1_a1_sumout),
	.datab(!fp_functions_0_aadd_1_a26_sumout),
	.datac(!fp_functions_0_aMux_59_a0_combout),
	.datad(!fp_functions_0_aMux_59_a1_combout),
	.datae(!fp_functions_0_aMux_59_a2_combout),
	.dataf(!fp_functions_0_aMux_59_a3_combout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai1783_a12_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai1783_a12.extended_lut = "off";
defparam fp_functions_0_ai1783_a12.lut_mask = 64'h02468ACE3377BBFF;
defparam fp_functions_0_ai1783_a12.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai1783_a13(
	.dataa(!fp_functions_0_aadd_1_a1_sumout),
	.datab(!fp_functions_0_aadd_1_a26_sumout),
	.datac(!fp_functions_0_aMux_60_a3_combout),
	.datad(!fp_functions_0_aMux_60_a4_combout),
	.datae(!fp_functions_0_aMux_76_a0_combout),
	.dataf(!fp_functions_0_aMux_60_a5_combout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai1783_a13_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai1783_a13.extended_lut = "off";
defparam fp_functions_0_ai1783_a13.lut_mask = 64'h0246CECE3377FFFF;
defparam fp_functions_0_ai1783_a13.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai1783_a14(
	.dataa(!fp_functions_0_aadd_1_a1_sumout),
	.datab(!fp_functions_0_aadd_1_a26_sumout),
	.datac(!fp_functions_0_aMux_59_a4_combout),
	.datad(!fp_functions_0_aMux_59_a5_combout),
	.datae(!fp_functions_0_aMux_59_a6_combout),
	.dataf(!fp_functions_0_aMux_79_a0_combout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai1783_a14_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai1783_a14.extended_lut = "off";
defparam fp_functions_0_ai1783_a14.lut_mask = 64'h01234567CDEFCDEF;
defparam fp_functions_0_ai1783_a14.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai1783_a15(
	.dataa(!fp_functions_0_aadd_1_a1_sumout),
	.datab(!fp_functions_0_aadd_1_a26_sumout),
	.datac(!fp_functions_0_aMux_58_a0_combout),
	.datad(!fp_functions_0_aMux_58_a1_combout),
	.datae(!fp_functions_0_aMux_78_a0_combout),
	.dataf(!fp_functions_0_aMux_62_a0_combout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai1783_a15_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai1783_a15.extended_lut = "off";
defparam fp_functions_0_ai1783_a15.lut_mask = 64'h0246CECE3377FFFF;
defparam fp_functions_0_ai1783_a15.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_50_a0(
	.dataa(!fp_functions_0_aadd_1_a16_sumout),
	.datab(!fp_functions_0_aadd_1_a21_sumout),
	.datac(!fp_functions_0_aadd_1_a1_sumout),
	.datad(!fp_functions_0_aMux_2_a20_combout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_50_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_50_a0.extended_lut = "off";
defparam fp_functions_0_aMux_50_a0.lut_mask = 64'h8000800080008000;
defparam fp_functions_0_aMux_50_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai1783_a16(
	.dataa(!fp_functions_0_aMux_58_a2_combout),
	.datab(!fp_functions_0_aMux_58_a3_combout),
	.datac(!fp_functions_0_aadd_1_a6_sumout),
	.datad(!fp_functions_0_aadd_3_a1_sumout),
	.datae(!fp_functions_0_ai1783_a32_combout),
	.dataf(!fp_functions_0_ai1783_a33_combout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai1783_a16_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai1783_a16.extended_lut = "off";
defparam fp_functions_0_ai1783_a16.lut_mask = 64'h000000F500000003;
defparam fp_functions_0_ai1783_a16.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_51_a0(
	.dataa(!fp_functions_0_afrac_bSig_uid36_fpAddTest_b_a21_a_a17_combout),
	.datab(!fp_functions_0_aadd_1_a16_sumout),
	.datac(!fp_functions_0_aadd_1_a21_sumout),
	.datad(!fp_functions_0_aadd_1_a1_sumout),
	.datae(!fp_functions_0_aMux_2_a11_combout),
	.dataf(!fp_functions_0_aMux_2_a12_combout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_51_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_51_a0.extended_lut = "off";
defparam fp_functions_0_aMux_51_a0.lut_mask = 64'h00007000C000F000;
defparam fp_functions_0_aMux_51_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai1783_a17(
	.dataa(!fp_functions_0_aadd_1_a1_sumout),
	.datab(!fp_functions_0_aMux_59_a0_combout),
	.datac(!fp_functions_0_aMux_59_a1_combout),
	.datad(!fp_functions_0_aadd_1_a6_sumout),
	.datae(!fp_functions_0_aadd_3_a1_sumout),
	.dataf(!fp_functions_0_ai1783_a30_combout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai1783_a17_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai1783_a17.extended_lut = "off";
defparam fp_functions_0_ai1783_a17.lut_mask = 64'h000000000000FF1B;
defparam fp_functions_0_ai1783_a17.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_52_a0(
	.dataa(!fp_functions_0_aadd_1_a16_sumout),
	.datab(!fp_functions_0_aadd_1_a21_sumout),
	.datac(!fp_functions_0_aMux_2_a17_combout),
	.datad(!fp_functions_0_aadd_1_a1_sumout),
	.datae(!fp_functions_0_areduce_nor_0_acombout),
	.dataf(!fp_functions_0_aMux_2_a20_combout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_52_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_52_a0.extended_lut = "off";
defparam fp_functions_0_aMux_52_a0.lut_mask = 64'h44004C0000000800;
defparam fp_functions_0_aMux_52_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai1783_a18(
	.dataa(!fp_functions_0_aadd_1_a1_sumout),
	.datab(!fp_functions_0_aMux_60_a3_combout),
	.datac(!fp_functions_0_aMux_60_a4_combout),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai1783_a18_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai1783_a18.extended_lut = "off";
defparam fp_functions_0_ai1783_a18.lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam fp_functions_0_ai1783_a18.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a13_a_a2(
	.dataa(!areset),
	.datab(!fp_functions_0_aadd_1_a21_sumout),
	.datac(!fp_functions_0_aadd_1_a1_sumout),
	.datad(!fp_functions_0_aadd_1_a6_sumout),
	.datae(!fp_functions_0_aadd_1_a26_sumout),
	.dataf(!fp_functions_0_aadd_3_a1_sumout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a13_a_a2_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a13_a_a2.extended_lut = "off";
defparam fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a13_a_a2.lut_mask = 64'hFFFFFFFFFDFF55FF;
defparam fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a13_a_a2.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai1783_a19(
	.dataa(!fp_functions_0_aadd_1_a1_sumout),
	.datab(!fp_functions_0_aMux_57_a3_combout),
	.datac(!fp_functions_0_aMux_57_a4_combout),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai1783_a19_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai1783_a19.extended_lut = "off";
defparam fp_functions_0_ai1783_a19.lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam fp_functions_0_ai1783_a19.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_53_a1(
	.dataa(!fp_functions_0_aadd_1_a16_sumout),
	.datab(!fp_functions_0_aadd_1_a21_sumout),
	.datac(!fp_functions_0_aadd_1_a1_sumout),
	.datad(!fp_functions_0_aMux_2_a11_combout),
	.datae(!fp_functions_0_aMux_2_a3_combout),
	.dataf(!fp_functions_0_aMux_2_a13_combout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_53_a1_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_53_a1.extended_lut = "off";
defparam fp_functions_0_aMux_53_a1.lut_mask = 64'h002080A04060C0E0;
defparam fp_functions_0_aMux_53_a1.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_54_a1(
	.dataa(!fp_functions_0_aadd_1_a16_sumout),
	.datab(!fp_functions_0_aadd_1_a21_sumout),
	.datac(!fp_functions_0_aadd_1_a1_sumout),
	.datad(!fp_functions_0_aMux_2_a19_combout),
	.datae(!fp_functions_0_aMux_2_a20_combout),
	.dataf(!fp_functions_0_aMux_2_a18_combout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_54_a1_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_54_a1.extended_lut = "off";
defparam fp_functions_0_aMux_54_a1.lut_mask = 64'h20A0008060E040C0;
defparam fp_functions_0_aMux_54_a1.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aexp_bSig_uid35_fpAddTest_b_a3_a_a0(
	.dataa(!b[26]),
	.datab(!a[26]),
	.datac(!fp_functions_0_aadd_0_a1_sumout),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aexp_bSig_uid35_fpAddTest_b_a3_a_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aexp_bSig_uid35_fpAddTest_b_a3_a_a0.extended_lut = "off";
defparam fp_functions_0_aexp_bSig_uid35_fpAddTest_b_a3_a_a0.lut_mask = 64'h5353535353535353;
defparam fp_functions_0_aexp_bSig_uid35_fpAddTest_b_a3_a_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aexp_bSig_uid35_fpAddTest_b_a1_a_a1(
	.dataa(!b[24]),
	.datab(!a[24]),
	.datac(!fp_functions_0_aadd_0_a1_sumout),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aexp_bSig_uid35_fpAddTest_b_a1_a_a1_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aexp_bSig_uid35_fpAddTest_b_a1_a_a1.extended_lut = "off";
defparam fp_functions_0_aexp_bSig_uid35_fpAddTest_b_a1_a_a1.lut_mask = 64'h5353535353535353;
defparam fp_functions_0_aexp_bSig_uid35_fpAddTest_b_a1_a_a1.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_areduce_nor_7_a0(
	.dataa(!b[23]),
	.datab(!a[23]),
	.datac(!fp_functions_0_aadd_0_a1_sumout),
	.datad(!fp_functions_0_aexp_bSig_uid35_fpAddTest_b_a1_a_a1_combout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_areduce_nor_7_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_areduce_nor_7_a0.extended_lut = "off";
defparam fp_functions_0_areduce_nor_7_a0.lut_mask = 64'hFFACFFACFFACFFAC;
defparam fp_functions_0_areduce_nor_7_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aexp_bSig_uid35_fpAddTest_b_a5_a_a2(
	.dataa(!b[28]),
	.datab(!a[28]),
	.datac(!fp_functions_0_aadd_0_a1_sumout),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aexp_bSig_uid35_fpAddTest_b_a5_a_a2_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aexp_bSig_uid35_fpAddTest_b_a5_a_a2.extended_lut = "off";
defparam fp_functions_0_aexp_bSig_uid35_fpAddTest_b_a5_a_a2.lut_mask = 64'h5353535353535353;
defparam fp_functions_0_aexp_bSig_uid35_fpAddTest_b_a5_a_a2.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_areduce_nor_7_a1(
	.dataa(!b[27]),
	.datab(!a[27]),
	.datac(!fp_functions_0_aadd_0_a1_sumout),
	.datad(!fp_functions_0_aexp_bSig_uid35_fpAddTest_b_a5_a_a2_combout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_areduce_nor_7_a1_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_areduce_nor_7_a1.extended_lut = "off";
defparam fp_functions_0_areduce_nor_7_a1.lut_mask = 64'hFFACFFACFFACFFAC;
defparam fp_functions_0_areduce_nor_7_a1.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aexp_bSig_uid35_fpAddTest_b_a7_a_a3(
	.dataa(!b[30]),
	.datab(!a[30]),
	.datac(!fp_functions_0_aadd_0_a1_sumout),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aexp_bSig_uid35_fpAddTest_b_a7_a_a3_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aexp_bSig_uid35_fpAddTest_b_a7_a_a3.extended_lut = "off";
defparam fp_functions_0_aexp_bSig_uid35_fpAddTest_b_a7_a_a3.lut_mask = 64'h5353535353535353;
defparam fp_functions_0_aexp_bSig_uid35_fpAddTest_b_a7_a_a3.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_areduce_nor_7_a2(
	.dataa(!b[29]),
	.datab(!a[29]),
	.datac(!fp_functions_0_aadd_0_a1_sumout),
	.datad(!fp_functions_0_aexp_bSig_uid35_fpAddTest_b_a7_a_a3_combout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_areduce_nor_7_a2_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_areduce_nor_7_a2.extended_lut = "off";
defparam fp_functions_0_areduce_nor_7_a2.lut_mask = 64'hFFACFFACFFACFFAC;
defparam fp_functions_0_areduce_nor_7_a2.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aexp_aSig_uid21_fpAddTest_b_a0_a_a0(
	.dataa(!b[27]),
	.datab(!a[27]),
	.datac(!fp_functions_0_aadd_0_a1_sumout),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aexp_aSig_uid21_fpAddTest_b_a0_a_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aexp_aSig_uid21_fpAddTest_b_a0_a_a0.extended_lut = "off";
defparam fp_functions_0_aexp_aSig_uid21_fpAddTest_b_a0_a_a0.lut_mask = 64'h3535353535353535;
defparam fp_functions_0_aexp_aSig_uid21_fpAddTest_b_a0_a_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aexp_aSig_uid21_fpAddTest_b_a0_a_a1(
	.dataa(!b[28]),
	.datab(!a[28]),
	.datac(!fp_functions_0_aadd_0_a1_sumout),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aexp_aSig_uid21_fpAddTest_b_a0_a_a1_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aexp_aSig_uid21_fpAddTest_b_a0_a_a1.extended_lut = "off";
defparam fp_functions_0_aexp_aSig_uid21_fpAddTest_b_a0_a_a1.lut_mask = 64'h3535353535353535;
defparam fp_functions_0_aexp_aSig_uid21_fpAddTest_b_a0_a_a1.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aexp_aSig_uid21_fpAddTest_b_a0_a_a2(
	.dataa(!b[29]),
	.datab(!a[29]),
	.datac(!fp_functions_0_aadd_0_a1_sumout),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aexp_aSig_uid21_fpAddTest_b_a0_a_a2_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aexp_aSig_uid21_fpAddTest_b_a0_a_a2.extended_lut = "off";
defparam fp_functions_0_aexp_aSig_uid21_fpAddTest_b_a0_a_a2.lut_mask = 64'h3535353535353535;
defparam fp_functions_0_aexp_aSig_uid21_fpAddTest_b_a0_a_a2.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aexp_aSig_uid21_fpAddTest_b_a0_a_a3(
	.dataa(!b[30]),
	.datab(!a[30]),
	.datac(!fp_functions_0_aadd_0_a1_sumout),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aexp_aSig_uid21_fpAddTest_b_a0_a_a3_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aexp_aSig_uid21_fpAddTest_b_a0_a_a3.extended_lut = "off";
defparam fp_functions_0_aexp_aSig_uid21_fpAddTest_b_a0_a_a3.lut_mask = 64'h3535353535353535;
defparam fp_functions_0_aexp_aSig_uid21_fpAddTest_b_a0_a_a3.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aexp_aSig_uid21_fpAddTest_b_a0_a_a4(
	.dataa(!b[23]),
	.datab(!a[23]),
	.datac(!fp_functions_0_aadd_0_a1_sumout),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aexp_aSig_uid21_fpAddTest_b_a0_a_a4_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aexp_aSig_uid21_fpAddTest_b_a0_a_a4.extended_lut = "off";
defparam fp_functions_0_aexp_aSig_uid21_fpAddTest_b_a0_a_a4.lut_mask = 64'h3535353535353535;
defparam fp_functions_0_aexp_aSig_uid21_fpAddTest_b_a0_a_a4.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aexp_aSig_uid21_fpAddTest_b_a0_a_a5(
	.dataa(!b[24]),
	.datab(!a[24]),
	.datac(!fp_functions_0_aadd_0_a1_sumout),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aexp_aSig_uid21_fpAddTest_b_a0_a_a5_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aexp_aSig_uid21_fpAddTest_b_a0_a_a5.extended_lut = "off";
defparam fp_functions_0_aexp_aSig_uid21_fpAddTest_b_a0_a_a5.lut_mask = 64'h3535353535353535;
defparam fp_functions_0_aexp_aSig_uid21_fpAddTest_b_a0_a_a5.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aexp_aSig_uid21_fpAddTest_b_a0_a_a6(
	.dataa(!b[25]),
	.datab(!a[25]),
	.datac(!fp_functions_0_aadd_0_a1_sumout),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aexp_aSig_uid21_fpAddTest_b_a0_a_a6_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aexp_aSig_uid21_fpAddTest_b_a0_a_a6.extended_lut = "off";
defparam fp_functions_0_aexp_aSig_uid21_fpAddTest_b_a0_a_a6.lut_mask = 64'h3535353535353535;
defparam fp_functions_0_aexp_aSig_uid21_fpAddTest_b_a0_a_a6.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aexp_aSig_uid21_fpAddTest_b_a0_a_a7(
	.dataa(!b[26]),
	.datab(!a[26]),
	.datac(!fp_functions_0_aadd_0_a1_sumout),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aexp_aSig_uid21_fpAddTest_b_a0_a_a7_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aexp_aSig_uid21_fpAddTest_b_a0_a_a7.extended_lut = "off";
defparam fp_functions_0_aexp_aSig_uid21_fpAddTest_b_a0_a_a7.lut_mask = 64'h3535353535353535;
defparam fp_functions_0_aexp_aSig_uid21_fpAddTest_b_a0_a_a7.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai326_a0(
	.dataa(!b[31]),
	.datab(!a[31]),
	.datac(!fp_functions_0_aadd_0_a1_sumout),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai326_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai326_a0.extended_lut = "off";
defparam fp_functions_0_ai326_a0.lut_mask = 64'h3535353535353535;
defparam fp_functions_0_ai326_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai289_a0(
	.dataa(!b[31]),
	.datab(!a[31]),
	.datac(!fp_functions_0_aadd_0_a1_sumout),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai289_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai289_a0.extended_lut = "off";
defparam fp_functions_0_ai289_a0.lut_mask = 64'h5353535353535353;
defparam fp_functions_0_ai289_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai2131_a0(
	.dataa(!b[19]),
	.datab(!a[19]),
	.datac(!fp_functions_0_aadd_0_a1_sumout),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai2131_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai2131_a0.extended_lut = "off";
defparam fp_functions_0_ai2131_a0.lut_mask = 64'h3535353535353535;
defparam fp_functions_0_ai2131_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai2131_a1(
	.dataa(!b[21]),
	.datab(!a[21]),
	.datac(!fp_functions_0_aadd_0_a1_sumout),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai2131_a1_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai2131_a1.extended_lut = "off";
defparam fp_functions_0_ai2131_a1.lut_mask = 64'h3535353535353535;
defparam fp_functions_0_ai2131_a1.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai2131_a2(
	.dataa(!b[15]),
	.datab(!a[15]),
	.datac(!fp_functions_0_aadd_0_a1_sumout),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai2131_a2_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai2131_a2.extended_lut = "off";
defparam fp_functions_0_ai2131_a2.lut_mask = 64'h3535353535353535;
defparam fp_functions_0_ai2131_a2.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai2131_a3(
	.dataa(!b[16]),
	.datab(!a[16]),
	.datac(!fp_functions_0_aadd_0_a1_sumout),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai2131_a3_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai2131_a3.extended_lut = "off";
defparam fp_functions_0_ai2131_a3.lut_mask = 64'h3535353535353535;
defparam fp_functions_0_ai2131_a3.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai2131_a4(
	.dataa(!b[17]),
	.datab(!a[17]),
	.datac(!fp_functions_0_aadd_0_a1_sumout),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai2131_a4_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai2131_a4.extended_lut = "off";
defparam fp_functions_0_ai2131_a4.lut_mask = 64'h3535353535353535;
defparam fp_functions_0_ai2131_a4.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai2131_a5(
	.dataa(!b[18]),
	.datab(!a[18]),
	.datac(!fp_functions_0_aadd_0_a1_sumout),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai2131_a5_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai2131_a5.extended_lut = "off";
defparam fp_functions_0_ai2131_a5.lut_mask = 64'h3535353535353535;
defparam fp_functions_0_ai2131_a5.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai2131_a6(
	.dataa(!b[20]),
	.datab(!a[20]),
	.datac(!fp_functions_0_aadd_0_a1_sumout),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai2131_a6_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai2131_a6.extended_lut = "off";
defparam fp_functions_0_ai2131_a6.lut_mask = 64'h3535353535353535;
defparam fp_functions_0_ai2131_a6.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai2131_a7(
	.dataa(!b[22]),
	.datab(!a[22]),
	.datac(!fp_functions_0_aadd_0_a1_sumout),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai2131_a7_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai2131_a7.extended_lut = "off";
defparam fp_functions_0_ai2131_a7.lut_mask = 64'h3535353535353535;
defparam fp_functions_0_ai2131_a7.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai2131_a8(
	.dataa(!b[2]),
	.datab(!a[2]),
	.datac(!fp_functions_0_aadd_0_a1_sumout),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai2131_a8_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai2131_a8.extended_lut = "off";
defparam fp_functions_0_ai2131_a8.lut_mask = 64'h3535353535353535;
defparam fp_functions_0_ai2131_a8.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai2131_a9(
	.dataa(!b[0]),
	.datab(!a[0]),
	.datac(!fp_functions_0_aadd_0_a1_sumout),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai2131_a9_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai2131_a9.extended_lut = "off";
defparam fp_functions_0_ai2131_a9.lut_mask = 64'h3535353535353535;
defparam fp_functions_0_ai2131_a9.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai2131_a10(
	.dataa(!b[1]),
	.datab(!a[1]),
	.datac(!fp_functions_0_aadd_0_a1_sumout),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai2131_a10_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai2131_a10.extended_lut = "off";
defparam fp_functions_0_ai2131_a10.lut_mask = 64'h3535353535353535;
defparam fp_functions_0_ai2131_a10.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai2131_a11(
	.dataa(!b[8]),
	.datab(!a[8]),
	.datac(!fp_functions_0_aadd_0_a1_sumout),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai2131_a11_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai2131_a11.extended_lut = "off";
defparam fp_functions_0_ai2131_a11.lut_mask = 64'h3535353535353535;
defparam fp_functions_0_ai2131_a11.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai2131_a12(
	.dataa(!b[13]),
	.datab(!a[13]),
	.datac(!fp_functions_0_aadd_0_a1_sumout),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai2131_a12_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai2131_a12.extended_lut = "off";
defparam fp_functions_0_ai2131_a12.lut_mask = 64'h3535353535353535;
defparam fp_functions_0_ai2131_a12.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai2131_a13(
	.dataa(!b[14]),
	.datab(!a[14]),
	.datac(!fp_functions_0_aadd_0_a1_sumout),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai2131_a13_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai2131_a13.extended_lut = "off";
defparam fp_functions_0_ai2131_a13.lut_mask = 64'h3535353535353535;
defparam fp_functions_0_ai2131_a13.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai2131_a14(
	.dataa(!b[9]),
	.datab(!a[9]),
	.datac(!fp_functions_0_aadd_0_a1_sumout),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai2131_a14_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai2131_a14.extended_lut = "off";
defparam fp_functions_0_ai2131_a14.lut_mask = 64'h3535353535353535;
defparam fp_functions_0_ai2131_a14.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai2131_a15(
	.dataa(!b[10]),
	.datab(!a[10]),
	.datac(!fp_functions_0_aadd_0_a1_sumout),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai2131_a15_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai2131_a15.extended_lut = "off";
defparam fp_functions_0_ai2131_a15.lut_mask = 64'h3535353535353535;
defparam fp_functions_0_ai2131_a15.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai2131_a16(
	.dataa(!b[11]),
	.datab(!a[11]),
	.datac(!fp_functions_0_aadd_0_a1_sumout),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai2131_a16_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai2131_a16.extended_lut = "off";
defparam fp_functions_0_ai2131_a16.lut_mask = 64'h3535353535353535;
defparam fp_functions_0_ai2131_a16.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai2131_a17(
	.dataa(!b[12]),
	.datab(!a[12]),
	.datac(!fp_functions_0_aadd_0_a1_sumout),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai2131_a17_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai2131_a17.extended_lut = "off";
defparam fp_functions_0_ai2131_a17.lut_mask = 64'h3535353535353535;
defparam fp_functions_0_ai2131_a17.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai2131_a18(
	.dataa(!b[3]),
	.datab(!a[3]),
	.datac(!fp_functions_0_aadd_0_a1_sumout),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai2131_a18_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai2131_a18.extended_lut = "off";
defparam fp_functions_0_ai2131_a18.lut_mask = 64'h3535353535353535;
defparam fp_functions_0_ai2131_a18.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai2131_a19(
	.dataa(!b[4]),
	.datab(!a[4]),
	.datac(!fp_functions_0_aadd_0_a1_sumout),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai2131_a19_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai2131_a19.extended_lut = "off";
defparam fp_functions_0_ai2131_a19.lut_mask = 64'h3535353535353535;
defparam fp_functions_0_ai2131_a19.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai2131_a20(
	.dataa(!b[5]),
	.datab(!a[5]),
	.datac(!fp_functions_0_aadd_0_a1_sumout),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai2131_a20_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai2131_a20.extended_lut = "off";
defparam fp_functions_0_ai2131_a20.lut_mask = 64'h3535353535353535;
defparam fp_functions_0_ai2131_a20.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai2131_a21(
	.dataa(!b[6]),
	.datab(!a[6]),
	.datac(!fp_functions_0_aadd_0_a1_sumout),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai2131_a21_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai2131_a21.extended_lut = "off";
defparam fp_functions_0_ai2131_a21.lut_mask = 64'h3535353535353535;
defparam fp_functions_0_ai2131_a21.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai2131_a22(
	.dataa(!b[7]),
	.datab(!a[7]),
	.datac(!fp_functions_0_aadd_0_a1_sumout),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai2131_a22_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai2131_a22.extended_lut = "off";
defparam fp_functions_0_ai2131_a22.lut_mask = 64'h3535353535353535;
defparam fp_functions_0_ai2131_a22.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_areduce_nor_10_a0(
	.dataa(!b[4]),
	.datab(!a[4]),
	.datac(!fp_functions_0_aadd_0_a1_sumout),
	.datad(!fp_functions_0_afrac_bSig_uid36_fpAddTest_b_a5_a_a8_combout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_areduce_nor_10_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_areduce_nor_10_a0.extended_lut = "off";
defparam fp_functions_0_areduce_nor_10_a0.lut_mask = 64'hAC00AC00AC00AC00;
defparam fp_functions_0_areduce_nor_10_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_areduce_nor_10_a1(
	.dataa(!b[1]),
	.datab(!a[1]),
	.datac(!b[0]),
	.datad(!a[0]),
	.datae(!fp_functions_0_aadd_0_a1_sumout),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_areduce_nor_10_a1_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_areduce_nor_10_a1.extended_lut = "off";
defparam fp_functions_0_areduce_nor_10_a1.lut_mask = 64'hA0A0CC00A0A0CC00;
defparam fp_functions_0_areduce_nor_10_a1.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_areduce_nor_10_a2(
	.dataa(!b[3]),
	.datab(!a[3]),
	.datac(!b[2]),
	.datad(!a[2]),
	.datae(!fp_functions_0_aadd_0_a1_sumout),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_areduce_nor_10_a2_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_areduce_nor_10_a2.extended_lut = "off";
defparam fp_functions_0_areduce_nor_10_a2.lut_mask = 64'hA0A0CC00A0A0CC00;
defparam fp_functions_0_areduce_nor_10_a2.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_areduce_nor_10_a3(
	.dataa(!fp_functions_0_afrac_bSig_uid36_fpAddTest_b_a19_a_a6_combout),
	.datab(!fp_functions_0_afrac_bSig_uid36_fpAddTest_b_a20_a_a7_combout),
	.datac(!fp_functions_0_afrac_bSig_uid36_fpAddTest_b_a21_a_a17_combout),
	.datad(!fp_functions_0_afrac_bSig_uid36_fpAddTest_b_a22_a_a18_combout),
	.datae(!fp_functions_0_areduce_nor_10_a1_combout),
	.dataf(!fp_functions_0_areduce_nor_10_a2_combout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_areduce_nor_10_a3_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_areduce_nor_10_a3.extended_lut = "off";
defparam fp_functions_0_areduce_nor_10_a3.lut_mask = 64'h0000000000008000;
defparam fp_functions_0_areduce_nor_10_a3.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_areduce_nor_10_a4(
	.dataa(!b[8]),
	.datab(!a[8]),
	.datac(!b[7]),
	.datad(!a[7]),
	.datae(!fp_functions_0_aadd_0_a1_sumout),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_areduce_nor_10_a4_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_areduce_nor_10_a4.extended_lut = "off";
defparam fp_functions_0_areduce_nor_10_a4.lut_mask = 64'hA0A0CC00A0A0CC00;
defparam fp_functions_0_areduce_nor_10_a4.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_areduce_nor_10_a5(
	.dataa(!b[12]),
	.datab(!a[12]),
	.datac(!b[11]),
	.datad(!a[11]),
	.datae(!fp_functions_0_aadd_0_a1_sumout),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_areduce_nor_10_a5_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_areduce_nor_10_a5.extended_lut = "off";
defparam fp_functions_0_areduce_nor_10_a5.lut_mask = 64'hA0A0CC00A0A0CC00;
defparam fp_functions_0_areduce_nor_10_a5.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_areduce_nor_10_a6(
	.dataa(!b[14]),
	.datab(!a[14]),
	.datac(!b[13]),
	.datad(!a[13]),
	.datae(!fp_functions_0_aadd_0_a1_sumout),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_areduce_nor_10_a6_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_areduce_nor_10_a6.extended_lut = "off";
defparam fp_functions_0_areduce_nor_10_a6.lut_mask = 64'hA0A0CC00A0A0CC00;
defparam fp_functions_0_areduce_nor_10_a6.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_areduce_nor_10_a7(
	.dataa(!b[16]),
	.datab(!a[16]),
	.datac(!b[15]),
	.datad(!a[15]),
	.datae(!fp_functions_0_aadd_0_a1_sumout),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_areduce_nor_10_a7_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_areduce_nor_10_a7.extended_lut = "off";
defparam fp_functions_0_areduce_nor_10_a7.lut_mask = 64'hA0A0CC00A0A0CC00;
defparam fp_functions_0_areduce_nor_10_a7.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_areduce_nor_10_a8(
	.dataa(!fp_functions_0_afrac_bSig_uid36_fpAddTest_b_a9_a_a12_combout),
	.datab(!fp_functions_0_afrac_bSig_uid36_fpAddTest_b_a10_a_a13_combout),
	.datac(!fp_functions_0_areduce_nor_10_a4_combout),
	.datad(!fp_functions_0_areduce_nor_10_a5_combout),
	.datae(!fp_functions_0_areduce_nor_10_a6_combout),
	.dataf(!fp_functions_0_areduce_nor_10_a7_combout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_areduce_nor_10_a8_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_areduce_nor_10_a8.extended_lut = "off";
defparam fp_functions_0_areduce_nor_10_a8.lut_mask = 64'h0000000000000008;
defparam fp_functions_0_areduce_nor_10_a8.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_areduce_nor_10(
	.dataa(!fp_functions_0_afrac_bSig_uid36_fpAddTest_b_a17_a_a4_combout),
	.datab(!fp_functions_0_afrac_bSig_uid36_fpAddTest_b_a18_a_a5_combout),
	.datac(!fp_functions_0_afrac_bSig_uid36_fpAddTest_b_a6_a_a9_combout),
	.datad(!fp_functions_0_areduce_nor_10_a0_combout),
	.datae(!fp_functions_0_areduce_nor_10_a3_combout),
	.dataf(!fp_functions_0_areduce_nor_10_a8_combout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_areduce_nor_10_acombout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_areduce_nor_10.extended_lut = "off";
defparam fp_functions_0_areduce_nor_10.lut_mask = 64'h0000000000000080;
defparam fp_functions_0_areduce_nor_10.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai3337_a3(
	.dataa(!fp_functions_0_areduce_nor_4_acombout),
	.datab(!fp_functions_0_arVStage_uid177_lzCountVal_uid85_fpAddTest_b_a0_a_a1_combout),
	.datac(!fp_functions_0_aMux_186_a1_combout),
	.datad(!fp_functions_0_aMux_186_a5_combout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai3337_a3_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai3337_a3.extended_lut = "off";
defparam fp_functions_0_ai3337_a3.lut_mask = 64'h0415041504150415;
defparam fp_functions_0_ai3337_a3.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai3337_a4(
	.dataa(!fp_functions_0_aredist1_vCount_uid152_lzCountVal_uid85_fpAddTest_q_1_q_a0_a_aq),
	.datab(!fp_functions_0_areduce_nor_3_acombout),
	.datac(!fp_functions_0_areduce_nor_6_a0_combout),
	.datad(!fp_functions_0_arVStage_uid165_lzCountVal_uid85_fpAddTest_merged_bit_select_b_a3_a_a6_combout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai3337_a4_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai3337_a4.extended_lut = "off";
defparam fp_functions_0_ai3337_a4.lut_mask = 64'h2220222022202220;
defparam fp_functions_0_ai3337_a4.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai3337_a5(
	.dataa(!fp_functions_0_aredist0_vStage_uid154_lzCountVal_uid85_fpAddTest_b_1_q_a1_a_aq),
	.datab(!fp_functions_0_ai3337_a4_combout),
	.datac(!fp_functions_0_areduce_nor_4_acombout),
	.datad(!fp_functions_0_arVStage_uid177_lzCountVal_uid85_fpAddTest_b_a0_a_a1_combout),
	.datae(!fp_functions_0_aMux_186_a5_combout),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai3337_a5_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai3337_a5.extended_lut = "off";
defparam fp_functions_0_ai3337_a5.lut_mask = 64'h00110F1100110F11;
defparam fp_functions_0_ai3337_a5.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai3337_a6(
	.dataa(!fp_functions_0_aredist0_vStage_uid154_lzCountVal_uid85_fpAddTest_b_1_q_a0_a_aq),
	.datab(!fp_functions_0_ai3337_a4_combout),
	.datac(!fp_functions_0_arVStage_uid177_lzCountVal_uid85_fpAddTest_b_a0_a_a1_combout),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai3337_a6_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai3337_a6.extended_lut = "off";
defparam fp_functions_0_ai3337_a6.lut_mask = 64'h1010101010101010;
defparam fp_functions_0_ai3337_a6.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai3337_a7(
	.dataa(!fp_functions_0_aredist0_vStage_uid154_lzCountVal_uid85_fpAddTest_b_1_q_a0_a_aq),
	.datab(!fp_functions_0_aredist0_vStage_uid154_lzCountVal_uid85_fpAddTest_b_1_q_a1_a_aq),
	.datac(!fp_functions_0_ai3337_a4_combout),
	.datad(!fp_functions_0_arVStage_uid177_lzCountVal_uid85_fpAddTest_b_a0_a_a1_combout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai3337_a7_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai3337_a7.extended_lut = "off";
defparam fp_functions_0_ai3337_a7.lut_mask = 64'h0305030503050305;
defparam fp_functions_0_ai3337_a7.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a41_a_a3(
	.dataa(!areset),
	.datab(!fp_functions_0_aadd_1_a6_sumout),
	.datac(!fp_functions_0_aadd_1_a26_sumout),
	.datad(!fp_functions_0_aadd_3_a1_sumout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a41_a_a3_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a41_a_a3.extended_lut = "off";
defparam fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a41_a_a3.lut_mask = 64'hFF7FFF7FFF7FFF7F;
defparam fp_functions_0_ar_uid219_alignmentShifter_uid64_fpAddTest_q_a41_a_a3.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_59_a7(
	.dataa(!fp_functions_0_aadd_1_a1_sumout),
	.datab(!fp_functions_0_aMux_59_a0_combout),
	.datac(!fp_functions_0_aMux_59_a3_combout),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_59_a7_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_59_a7.extended_lut = "off";
defparam fp_functions_0_aMux_59_a7.lut_mask = 64'h2F2F2F2F2F2F2F2F;
defparam fp_functions_0_aMux_59_a7.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_63_a0(
	.dataa(!fp_functions_0_aadd_1_a1_sumout),
	.datab(!fp_functions_0_aMux_59_a4_combout),
	.datac(!fp_functions_0_aMux_59_a5_combout),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_63_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_63_a0.extended_lut = "off";
defparam fp_functions_0_aMux_63_a0.lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam fp_functions_0_aMux_63_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_62_a1(
	.dataa(!fp_functions_0_aadd_1_a1_sumout),
	.datab(!fp_functions_0_aMux_58_a0_combout),
	.datac(!fp_functions_0_aMux_62_a0_combout),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_62_a1_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_62_a1.extended_lut = "off";
defparam fp_functions_0_aMux_62_a1.lut_mask = 64'h2F2F2F2F2F2F2F2F;
defparam fp_functions_0_aMux_62_a1.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_61_a1(
	.dataa(!fp_functions_0_aadd_1_a1_sumout),
	.datab(!fp_functions_0_aMux_57_a3_combout),
	.datac(!fp_functions_0_aMux_61_a0_combout),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_61_a1_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_61_a1.extended_lut = "off";
defparam fp_functions_0_aMux_61_a1.lut_mask = 64'h2F2F2F2F2F2F2F2F;
defparam fp_functions_0_aMux_61_a1.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_60_a6(
	.dataa(!fp_functions_0_aadd_1_a1_sumout),
	.datab(!fp_functions_0_aMux_60_a3_combout),
	.datac(!fp_functions_0_aMux_60_a5_combout),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_60_a6_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_60_a6.extended_lut = "off";
defparam fp_functions_0_aMux_60_a6.lut_mask = 64'h2F2F2F2F2F2F2F2F;
defparam fp_functions_0_aMux_60_a6.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_58_a5(
	.dataa(!fp_functions_0_aadd_1_a1_sumout),
	.datab(!fp_functions_0_aMux_58_a2_combout),
	.datac(!fp_functions_0_aMux_58_a4_combout),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_58_a5_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_58_a5.extended_lut = "off";
defparam fp_functions_0_aMux_58_a5.lut_mask = 64'h2F2F2F2F2F2F2F2F;
defparam fp_functions_0_aMux_58_a5.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_57_a6(
	.dataa(!fp_functions_0_aadd_1_a1_sumout),
	.datab(!fp_functions_0_aMux_57_a0_combout),
	.datac(!fp_functions_0_aMux_57_a5_combout),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_57_a6_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_57_a6.extended_lut = "off";
defparam fp_functions_0_aMux_57_a6.lut_mask = 64'h2F2F2F2F2F2F2F2F;
defparam fp_functions_0_aMux_57_a6.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_56_a1(
	.dataa(!fp_functions_0_aadd_1_a1_sumout),
	.datab(!fp_functions_0_aMux_60_a0_combout),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_56_a1_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_56_a1.extended_lut = "off";
defparam fp_functions_0_aMux_56_a1.lut_mask = 64'h2222222222222222;
defparam fp_functions_0_aMux_56_a1.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai1783_a20(
	.dataa(!fp_functions_0_aadd_1_a1_sumout),
	.datab(!fp_functions_0_aadd_1_a6_sumout),
	.datac(!fp_functions_0_aMux_60_a3_combout),
	.datad(!fp_functions_0_aMux_60_a4_combout),
	.datae(!fp_functions_0_aMux_52_a0_combout),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai1783_a20_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai1783_a20.extended_lut = "off";
defparam fp_functions_0_ai1783_a20.lut_mask = 64'h048C37BF048C37BF;
defparam fp_functions_0_ai1783_a20.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai1783_a21(
	.dataa(!fp_functions_0_aadd_1_a1_sumout),
	.datab(!fp_functions_0_aadd_1_a6_sumout),
	.datac(!fp_functions_0_aMux_57_a3_combout),
	.datad(!fp_functions_0_aMux_57_a4_combout),
	.datae(!fp_functions_0_aMux_53_a1_combout),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai1783_a21_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai1783_a21.extended_lut = "off";
defparam fp_functions_0_ai1783_a21.lut_mask = 64'h048C37BF048C37BF;
defparam fp_functions_0_ai1783_a21.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai1783_a22(
	.dataa(!fp_functions_0_aadd_1_a1_sumout),
	.datab(!fp_functions_0_aadd_1_a6_sumout),
	.datac(!fp_functions_0_aMux_59_a4_combout),
	.datad(!fp_functions_0_aMux_59_a5_combout),
	.datae(!fp_functions_0_aMux_59_a6_combout),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai1783_a22_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai1783_a22.extended_lut = "off";
defparam fp_functions_0_ai1783_a22.lut_mask = 64'h02468ACE02468ACE;
defparam fp_functions_0_ai1783_a22.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai1783_a23(
	.dataa(!fp_functions_0_aadd_1_a1_sumout),
	.datab(!fp_functions_0_aadd_1_a6_sumout),
	.datac(!fp_functions_0_aMux_58_a0_combout),
	.datad(!fp_functions_0_aMux_58_a1_combout),
	.datae(!fp_functions_0_aMux_54_a1_combout),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai1783_a23_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai1783_a23.extended_lut = "off";
defparam fp_functions_0_ai1783_a23.lut_mask = 64'h048C37BF048C37BF;
defparam fp_functions_0_ai1783_a23.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_aMux_64_a0(
	.dataa(!fp_functions_0_aadd_1_a1_sumout),
	.datab(!fp_functions_0_aMux_60_a0_combout),
	.datac(!fp_functions_0_aMux_60_a1_combout),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_aMux_64_a0_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_aMux_64_a0.extended_lut = "off";
defparam fp_functions_0_aMux_64_a0.lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam fp_functions_0_aMux_64_a0.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai1783_a24(
	.dataa(!fp_functions_0_aadd_1_a1_sumout),
	.datab(!fp_functions_0_aadd_1_a6_sumout),
	.datac(!fp_functions_0_aMux_57_a0_combout),
	.datad(!fp_functions_0_aMux_57_a1_combout),
	.datae(!fp_functions_0_aMux_49_a0_combout),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai1783_a24_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai1783_a24.extended_lut = "off";
defparam fp_functions_0_ai1783_a24.lut_mask = 64'h048C37BF048C37BF;
defparam fp_functions_0_ai1783_a24.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai1783_a25(
	.dataa(!fp_functions_0_aadd_1_a1_sumout),
	.datab(!fp_functions_0_aadd_1_a6_sumout),
	.datac(!fp_functions_0_aMux_60_a0_combout),
	.datad(!fp_functions_0_aMux_60_a1_combout),
	.datae(!fp_functions_0_aMux_60_a2_combout),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai1783_a25_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai1783_a25.extended_lut = "off";
defparam fp_functions_0_ai1783_a25.lut_mask = 64'h02468ACE02468ACE;
defparam fp_functions_0_ai1783_a25.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai1783_a26(
	.dataa(!fp_functions_0_aadd_1_a1_sumout),
	.datab(!fp_functions_0_aadd_1_a6_sumout),
	.datac(!fp_functions_0_aMux_59_a0_combout),
	.datad(!fp_functions_0_aMux_59_a1_combout),
	.datae(!fp_functions_0_aMux_51_a0_combout),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai1783_a26_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai1783_a26.extended_lut = "off";
defparam fp_functions_0_ai1783_a26.lut_mask = 64'h048C37BF048C37BF;
defparam fp_functions_0_ai1783_a26.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai1783_a27(
	.dataa(!fp_functions_0_aadd_1_a1_sumout),
	.datab(!fp_functions_0_aadd_1_a6_sumout),
	.datac(!fp_functions_0_aMux_58_a2_combout),
	.datad(!fp_functions_0_aMux_58_a3_combout),
	.datae(!fp_functions_0_aMux_50_a0_combout),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai1783_a27_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai1783_a27.extended_lut = "off";
defparam fp_functions_0_ai1783_a27.lut_mask = 64'h048C37BF048C37BF;
defparam fp_functions_0_ai1783_a27.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai1783_a28(
	.dataa(!fp_functions_0_aadd_1_a1_sumout),
	.datab(!fp_functions_0_aadd_1_a6_sumout),
	.datac(!fp_functions_0_aMux_57_a0_combout),
	.datad(!fp_functions_0_aMux_57_a1_combout),
	.datae(!fp_functions_0_aMux_57_a5_combout),
	.dataf(!fp_functions_0_aMux_57_a2_combout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai1783_a28_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai1783_a28.extended_lut = "off";
defparam fp_functions_0_ai1783_a28.lut_mask = 64'h024633778ACEBBFF;
defparam fp_functions_0_ai1783_a28.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai1783_a29(
	.dataa(!fp_functions_0_aadd_1_a1_sumout),
	.datab(!fp_functions_0_aadd_1_a6_sumout),
	.datac(!fp_functions_0_aMux_58_a2_combout),
	.datad(!fp_functions_0_aMux_58_a3_combout),
	.datae(!fp_functions_0_aMux_58_a4_combout),
	.dataf(!fp_functions_0_ai1783_a10_combout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai1783_a29_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai1783_a29.extended_lut = "off";
defparam fp_functions_0_ai1783_a29.lut_mask = 64'h02463377CECEFFFF;
defparam fp_functions_0_ai1783_a29.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai1783_a30(
	.dataa(!fp_functions_0_aMux_59_a2_combout),
	.datab(!fp_functions_0_aMux_51_a0_combout),
	.datac(!fp_functions_0_aadd_1_a1_sumout),
	.datad(!areset),
	.datae(!fp_functions_0_aadd_1_a6_sumout),
	.dataf(!fp_functions_0_aadd_1_a26_sumout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai1783_a30_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai1783_a30.extended_lut = "off";
defparam fp_functions_0_ai1783_a30.lut_mask = 64'h0500FF0033000000;
defparam fp_functions_0_ai1783_a30.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai1783_a31(
	.dataa(!fp_functions_0_aadd_1_a16_sumout),
	.datab(!fp_functions_0_aadd_1_a21_sumout),
	.datac(!fp_functions_0_aMux_23_a0_combout),
	.datad(!fp_functions_0_aMux_23_a1_combout),
	.datae(!fp_functions_0_aMux_2_a26_combout),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai1783_a31_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai1783_a31.extended_lut = "off";
defparam fp_functions_0_ai1783_a31.lut_mask = 64'h0426153704261537;
defparam fp_functions_0_ai1783_a31.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai1783_a32(
	.dataa(!fp_functions_0_aMux_50_a0_combout),
	.datab(!fp_functions_0_aadd_1_a1_sumout),
	.datac(!areset),
	.datad(!fp_functions_0_aadd_1_a6_sumout),
	.datae(!fp_functions_0_aadd_1_a26_sumout),
	.dataf(!fp_functions_0_areduce_nor_0_acombout),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai1783_a32_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai1783_a32.extended_lut = "off";
defparam fp_functions_0_ai1783_a32.lut_mask = 64'h00F0500030F05000;
defparam fp_functions_0_ai1783_a32.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_ai1783_a33(
	.dataa(!fp_functions_0_aadd_1_a1_sumout),
	.datab(!fp_functions_0_aadd_1_a6_sumout),
	.datac(!fp_functions_0_aadd_1_a26_sumout),
	.datad(!fp_functions_0_ai1783_a31_combout),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_ai1783_a33_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_ai1783_a33.extended_lut = "off";
defparam fp_functions_0_ai1783_a33.lut_mask = 64'hE0A0E0A0E0A0E0A0;
defparam fp_functions_0_ai1783_a33.shared_arith = "off";

fourteennm_lcell_comb fp_functions_0_areduce_nor_0_a_wirecell(
	.dataa(!fp_functions_0_areduce_nor_0_acombout),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fp_functions_0_areduce_nor_0_a_wirecell_combout),
	.sumout(),
	.cout(),
	.shareout());
defparam fp_functions_0_areduce_nor_0_a_wirecell.extended_lut = "off";
defparam fp_functions_0_areduce_nor_0_a_wirecell.lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam fp_functions_0_areduce_nor_0_a_wirecell.shared_arith = "off";

assign q[30] = fp_functions_0_aMux_207_a2_combout;

assign q[29] = fp_functions_0_aMux_208_a2_combout;

assign q[28] = fp_functions_0_aMux_209_a2_combout;

assign q[27] = fp_functions_0_aMux_210_a2_combout;

assign q[26] = fp_functions_0_aMux_211_a2_combout;

assign q[25] = fp_functions_0_aMux_212_a2_combout;

assign q[24] = fp_functions_0_aMux_213_a2_combout;

assign q[23] = fp_functions_0_aMux_214_a2_combout;

assign q[22] = fp_functions_0_aMux_215_a0_combout;

assign q[21] = fp_functions_0_aMux_216_a0_combout;

assign q[20] = fp_functions_0_aMux_217_a0_combout;

assign q[19] = fp_functions_0_aMux_218_a0_combout;

assign q[18] = fp_functions_0_aMux_219_a0_combout;

assign q[17] = fp_functions_0_aMux_220_a0_combout;

assign q[16] = fp_functions_0_aMux_221_a0_combout;

assign q[15] = fp_functions_0_aMux_222_a0_combout;

assign q[14] = fp_functions_0_aMux_223_a0_combout;

assign q[13] = fp_functions_0_aMux_224_a0_combout;

assign q[12] = fp_functions_0_aMux_225_a0_combout;

assign q[11] = fp_functions_0_aMux_226_a0_combout;

assign q[10] = fp_functions_0_aMux_227_a0_combout;

assign q[9] = fp_functions_0_aMux_228_a0_combout;

assign q[8] = fp_functions_0_aMux_229_a0_combout;

assign q[7] = fp_functions_0_aMux_230_a0_combout;

assign q[6] = fp_functions_0_aMux_231_a0_combout;

assign q[5] = fp_functions_0_aMux_232_a0_combout;

assign q[4] = fp_functions_0_aMux_233_a0_combout;

assign q[3] = fp_functions_0_aMux_234_a0_combout;

assign q[2] = fp_functions_0_aMux_235_a0_combout;

assign q[1] = fp_functions_0_aMux_236_a1_combout;

assign q[0] = fp_functions_0_aMux_237_a2_combout;

assign q[31] = fp_functions_0_aR_uid148_fpAddTest_q_a31_a_a0_combout;

endmodule
